VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO IMPACTSram
  CLASS BLOCK ;
  FOREIGN IMPACTSram ;
  ORIGIN 0.790 43.350 ;
  SIZE 221.940 BY 67.830 ;
  PIN BL0
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met1 ;
        RECT 1.660 18.680 1.680 18.700 ;
        RECT 1.300 -43.100 1.980 -41.550 ;
    END
  END BL0
  PIN BLb0
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met1 ;
        RECT 6.780 18.630 6.800 18.650 ;
        RECT 6.400 -43.120 7.080 -41.550 ;
    END
  END BLb0
  PIN BL1
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met1 ;
        RECT 8.390 18.590 8.410 18.610 ;
        RECT 8.040 -43.110 8.720 -41.550 ;
    END
  END BL1
  PIN BLb1
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met1 ;
        RECT 13.540 18.470 13.560 18.490 ;
        RECT 13.160 -43.110 13.840 -41.550 ;
    END
  END BLb1
  PIN BL2
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met1 ;
        RECT 15.150 18.510 15.170 18.530 ;
        RECT 14.800 -43.110 15.480 -41.550 ;
    END
  END BL2
  PIN BLb2
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met1 ;
        RECT 20.310 18.700 20.330 18.720 ;
        RECT 19.910 -43.120 20.590 -41.550 ;
    END
  END BLb2
  PIN BL3
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met1 ;
        RECT 21.870 18.620 21.890 18.640 ;
        RECT 21.550 -43.110 22.230 -41.550 ;
    END
  END BL3
  PIN BLb3
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met1 ;
        RECT 26.990 18.690 27.010 18.710 ;
        RECT 26.650 -43.100 27.330 -41.550 ;
    END
  END BLb3
  PIN BL4
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met1 ;
        RECT 28.690 18.720 28.710 18.740 ;
        RECT 28.300 -43.100 28.980 -41.550 ;
    END
  END BL4
  PIN BLb4
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met1 ;
        RECT 33.780 18.700 33.800 18.720 ;
        RECT 33.400 -43.110 34.080 -41.550 ;
    END
  END BLb4
  PIN BL5
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met1 ;
        RECT 35.450 18.690 35.470 18.710 ;
        RECT 35.040 -43.120 35.720 -41.550 ;
    END
  END BL5
  PIN BLb5
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met1 ;
        RECT 40.530 18.460 40.550 18.480 ;
        RECT 40.150 -43.110 40.830 -41.550 ;
    END
  END BLb5
  PIN BL6
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met1 ;
        RECT 42.170 18.510 42.190 18.530 ;
        RECT 41.790 -43.110 42.470 -41.550 ;
    END
  END BL6
  PIN BLb6
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met1 ;
        RECT 47.280 18.350 47.300 18.370 ;
        RECT 46.910 -43.110 47.590 -41.550 ;
    END
  END BLb6
  PIN BL7
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met1 ;
        RECT 48.930 18.780 48.950 18.800 ;
        RECT 48.550 -43.120 49.230 -41.550 ;
    END
  END BL7
  PIN BLb7
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met1 ;
        RECT 53.970 18.680 53.990 18.700 ;
        RECT 53.650 -43.100 54.330 -41.550 ;
    END
  END BLb7
  PIN BL8
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met1 ;
        RECT 55.680 18.700 55.700 18.720 ;
        RECT 55.300 -43.100 55.980 -41.550 ;
    END
  END BL8
  PIN BLb8
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met1 ;
        RECT 60.870 18.720 60.890 18.740 ;
        RECT 60.400 -43.120 61.080 -41.550 ;
    END
  END BLb8
  PIN BL9
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met1 ;
        RECT 62.410 18.820 62.430 18.840 ;
        RECT 62.040 -43.110 62.720 -41.550 ;
    END
  END BL9
  PIN BLb9
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met1 ;
        RECT 67.510 18.850 67.530 18.870 ;
        RECT 67.160 -43.110 67.840 -41.550 ;
    END
  END BLb9
  PIN BL10
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met1 ;
        RECT 69.120 18.820 69.140 18.840 ;
        RECT 68.800 -43.110 69.480 -41.550 ;
    END
  END BL10
  PIN BLb10
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met1 ;
        RECT 74.310 18.820 74.330 18.840 ;
        RECT 73.910 -43.120 74.590 -41.550 ;
    END
  END BLb10
  PIN BL11
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met1 ;
        RECT 75.910 18.810 75.930 18.830 ;
        RECT 75.550 -43.110 76.230 -41.550 ;
    END
  END BL11
  PIN BLb11
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met1 ;
        RECT 81.040 18.890 81.060 18.910 ;
        RECT 80.650 -43.100 81.330 -41.550 ;
    END
  END BLb11
  PIN BL12
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met1 ;
        RECT 82.640 18.620 82.660 18.640 ;
        RECT 82.300 -43.100 82.980 -41.550 ;
    END
  END BL12
  PIN BLb12
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met1 ;
        RECT 87.780 18.510 87.800 18.530 ;
        RECT 87.400 -43.110 88.080 -41.550 ;
    END
  END BLb12
  PIN BL13
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met1 ;
        RECT 89.410 18.560 89.430 18.580 ;
        RECT 89.040 -43.120 89.720 -41.550 ;
    END
  END BL13
  PIN BLb13
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met1 ;
        RECT 94.530 18.550 94.550 18.570 ;
        RECT 94.150 -43.110 94.830 -41.550 ;
    END
  END BLb13
  PIN BL14
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met1 ;
        RECT 96.150 18.390 96.170 18.410 ;
        RECT 95.790 -43.110 96.470 -41.550 ;
    END
  END BL14
  PIN BLb14
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met1 ;
        RECT 101.310 18.490 101.330 18.510 ;
        RECT 100.910 -43.110 101.590 -41.550 ;
    END
  END BLb14
  PIN BL15
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met1 ;
        RECT 102.870 18.600 102.890 18.620 ;
        RECT 102.550 -43.120 103.230 -41.550 ;
    END
  END BL15
  PIN BLb15
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met1 ;
        RECT 108.020 18.410 108.040 18.430 ;
        RECT 107.650 -43.100 108.330 -41.550 ;
    END
  END BLb15
  PIN WL0
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER li1 ;
        RECT 0.590 15.310 1.010 15.750 ;
      LAYER mcon ;
        RECT 0.680 15.400 0.950 15.670 ;
      LAYER met1 ;
        RECT 0.590 15.760 1.010 16.230 ;
        RECT 0.580 15.310 1.010 15.760 ;
      LAYER via ;
        RECT 0.680 15.900 0.950 16.170 ;
      LAYER met2 ;
        RECT 0.580 15.760 1.010 16.270 ;
        RECT 0.590 15.750 1.010 15.760 ;
    END
  END WL0
  PIN WL1
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER li1 ;
        RECT 0.590 14.420 1.010 14.860 ;
      LAYER mcon ;
        RECT 0.680 14.500 0.950 14.770 ;
      LAYER met1 ;
        RECT 0.580 14.410 1.010 14.860 ;
        RECT 0.590 13.940 1.010 14.410 ;
      LAYER via ;
        RECT 0.680 14.000 0.950 14.270 ;
      LAYER met2 ;
        RECT 0.590 13.900 1.010 14.430 ;
    END
  END WL1
  PIN WL2
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER li1 ;
        RECT 0.590 11.700 1.010 12.140 ;
      LAYER mcon ;
        RECT 0.680 11.790 0.950 12.060 ;
      LAYER met1 ;
        RECT 0.590 12.150 1.010 12.620 ;
        RECT 0.580 11.700 1.010 12.150 ;
      LAYER via ;
        RECT 0.680 12.290 0.950 12.560 ;
      LAYER met2 ;
        RECT 0.590 12.630 1.010 12.670 ;
        RECT 0.580 12.150 1.010 12.630 ;
        RECT 0.590 12.140 1.010 12.150 ;
    END
  END WL2
  PIN WL3
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER li1 ;
        RECT 0.590 10.810 1.010 11.250 ;
      LAYER mcon ;
        RECT 0.680 10.890 0.950 11.160 ;
      LAYER met1 ;
        RECT 0.580 10.800 1.010 11.250 ;
        RECT 0.590 10.330 1.010 10.800 ;
      LAYER via ;
        RECT 0.680 10.390 0.950 10.660 ;
      LAYER met2 ;
        RECT 0.590 10.790 1.010 10.820 ;
        RECT 0.580 10.310 1.010 10.790 ;
        RECT 1.040 10.460 1.060 10.480 ;
        RECT 0.590 10.300 1.010 10.310 ;
    END
  END WL3
  PIN WL4
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER li1 ;
        RECT 0.590 8.090 1.010 8.530 ;
      LAYER mcon ;
        RECT 0.680 8.180 0.950 8.450 ;
      LAYER met1 ;
        RECT 0.590 8.540 1.010 9.010 ;
        RECT 0.580 8.090 1.010 8.540 ;
      LAYER via ;
        RECT 0.680 8.680 0.950 8.950 ;
      LAYER met2 ;
        RECT 0.580 8.670 1.010 9.050 ;
        RECT 0.580 8.650 1.020 8.670 ;
        RECT 0.580 8.540 1.010 8.650 ;
        RECT 0.590 8.520 1.010 8.540 ;
    END
  END WL4
  PIN WL5
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER li1 ;
        RECT 0.590 7.200 1.010 7.640 ;
      LAYER mcon ;
        RECT 0.680 7.280 0.950 7.550 ;
      LAYER met1 ;
        RECT 0.580 7.190 1.010 7.640 ;
        RECT 0.590 6.720 1.010 7.190 ;
      LAYER via ;
        RECT 0.680 6.780 0.950 7.050 ;
      LAYER met2 ;
        RECT 0.880 7.200 1.010 7.210 ;
        RECT 0.590 7.190 1.010 7.200 ;
        RECT 0.580 6.670 1.010 7.190 ;
        RECT 1.020 7.100 1.040 7.120 ;
    END
  END WL5
  PIN WL6
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER li1 ;
        RECT 0.590 4.480 1.010 4.920 ;
      LAYER mcon ;
        RECT 0.680 4.570 0.950 4.840 ;
      LAYER met1 ;
        RECT 0.590 4.930 1.010 5.400 ;
        RECT 0.580 4.480 1.010 4.930 ;
      LAYER via ;
        RECT 0.680 5.070 0.950 5.340 ;
      LAYER met2 ;
        RECT 0.590 4.910 1.010 5.430 ;
        RECT 1.050 5.240 1.070 5.260 ;
    END
  END WL6
  PIN WL7
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER li1 ;
        RECT 0.590 3.590 1.010 4.030 ;
      LAYER mcon ;
        RECT 0.680 3.670 0.950 3.940 ;
      LAYER met1 ;
        RECT 0.580 3.580 1.010 4.030 ;
        RECT 0.590 3.110 1.010 3.580 ;
      LAYER via ;
        RECT 0.680 3.170 0.950 3.440 ;
      LAYER met2 ;
        RECT 0.590 3.570 1.010 3.590 ;
        RECT 0.580 3.490 1.010 3.570 ;
        RECT 0.580 3.470 1.030 3.490 ;
        RECT 0.580 3.060 1.010 3.470 ;
    END
  END WL7
  PIN WL8
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER li1 ;
        RECT 0.590 0.870 1.010 1.310 ;
      LAYER mcon ;
        RECT 0.680 0.960 0.950 1.230 ;
      LAYER met1 ;
        RECT 0.590 1.320 1.010 1.790 ;
        RECT 0.580 0.870 1.010 1.320 ;
      LAYER via ;
        RECT 0.680 1.460 0.950 1.730 ;
      LAYER met2 ;
        RECT 0.580 1.330 1.010 1.840 ;
        RECT 1.030 1.590 1.050 1.610 ;
        RECT 0.590 1.310 1.010 1.330 ;
    END
  END WL8
  PIN WL9
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER li1 ;
        RECT 0.590 -0.020 1.010 0.420 ;
      LAYER mcon ;
        RECT 0.680 0.060 0.950 0.330 ;
      LAYER met1 ;
        RECT 0.580 -0.030 1.010 0.420 ;
        RECT 0.590 -0.500 1.010 -0.030 ;
      LAYER via ;
        RECT 0.680 -0.440 0.950 -0.170 ;
      LAYER met2 ;
        RECT 0.590 -0.530 1.010 -0.010 ;
        RECT 1.050 -0.160 1.070 -0.140 ;
    END
  END WL9
  PIN WL10
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER li1 ;
        RECT 0.590 -2.740 1.010 -2.300 ;
      LAYER mcon ;
        RECT 0.680 -2.650 0.950 -2.380 ;
      LAYER met1 ;
        RECT 0.590 -2.290 1.010 -1.820 ;
        RECT 0.580 -2.740 1.010 -2.290 ;
      LAYER via ;
        RECT 0.680 -2.150 0.950 -1.880 ;
      LAYER met2 ;
        RECT 0.580 -2.290 1.010 -1.770 ;
        RECT 1.030 -1.870 1.050 -1.850 ;
        RECT 0.590 -2.300 1.010 -2.290 ;
    END
  END WL10
  PIN WL11
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER li1 ;
        RECT 0.590 -3.630 1.010 -3.190 ;
      LAYER mcon ;
        RECT 0.680 -3.550 0.950 -3.280 ;
      LAYER met1 ;
        RECT 0.580 -3.640 1.010 -3.190 ;
        RECT 0.590 -4.110 1.010 -3.640 ;
      LAYER via ;
        RECT 0.680 -4.050 0.950 -3.780 ;
      LAYER met2 ;
        RECT 0.590 -3.640 1.010 -3.620 ;
        RECT 0.580 -4.150 1.010 -3.640 ;
        RECT 1.020 -3.710 1.040 -3.690 ;
    END
  END WL11
  PIN WL12
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER li1 ;
        RECT 0.590 -6.350 1.010 -5.910 ;
      LAYER mcon ;
        RECT 0.680 -6.260 0.950 -5.990 ;
      LAYER met1 ;
        RECT 0.590 -5.900 1.010 -5.430 ;
        RECT 0.580 -6.350 1.010 -5.900 ;
      LAYER via ;
        RECT 0.680 -5.760 0.950 -5.490 ;
      LAYER met2 ;
        RECT 0.870 -5.400 1.010 -5.390 ;
        RECT 0.590 -5.410 1.010 -5.400 ;
        RECT 0.580 -5.460 1.010 -5.410 ;
        RECT 0.580 -5.480 1.030 -5.460 ;
        RECT 0.580 -5.890 1.010 -5.480 ;
        RECT 0.590 -5.920 1.010 -5.890 ;
    END
  END WL12
  PIN WL13
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER li1 ;
        RECT 0.590 -7.240 1.010 -6.800 ;
      LAYER mcon ;
        RECT 0.680 -7.160 0.950 -6.890 ;
      LAYER met1 ;
        RECT 0.580 -7.250 1.010 -6.800 ;
        RECT 0.590 -7.720 1.010 -7.250 ;
      LAYER via ;
        RECT 0.680 -7.660 0.950 -7.390 ;
      LAYER met2 ;
        RECT 0.590 -7.250 1.010 -7.240 ;
        RECT 0.580 -7.730 1.010 -7.250 ;
        RECT 1.030 -7.550 1.050 -7.530 ;
        RECT 0.590 -7.770 1.010 -7.730 ;
    END
  END WL13
  PIN WL14
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER li1 ;
        RECT 0.590 -9.960 1.010 -9.520 ;
      LAYER mcon ;
        RECT 0.680 -9.870 0.950 -9.600 ;
      LAYER met1 ;
        RECT 0.590 -9.510 1.010 -9.040 ;
        RECT 0.580 -9.960 1.010 -9.510 ;
      LAYER via ;
        RECT 0.680 -9.370 0.950 -9.100 ;
      LAYER met2 ;
        RECT 0.590 -9.240 1.010 -9.000 ;
        RECT 0.590 -9.260 1.030 -9.240 ;
        RECT 0.590 -9.530 1.010 -9.260 ;
    END
  END WL14
  PIN WL15
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER li1 ;
        RECT 0.590 -10.850 1.010 -10.410 ;
      LAYER mcon ;
        RECT 0.680 -10.770 0.950 -10.500 ;
      LAYER met1 ;
        RECT 0.580 -10.860 1.010 -10.410 ;
        RECT 0.590 -11.330 1.010 -10.860 ;
      LAYER via ;
        RECT 0.680 -11.270 0.950 -11.000 ;
      LAYER met2 ;
        RECT 0.590 -10.860 1.010 -10.850 ;
        RECT 0.580 -10.950 1.010 -10.860 ;
        RECT 0.580 -10.970 1.030 -10.950 ;
        RECT 0.580 -11.370 1.010 -10.970 ;
    END
  END WL15
  PIN WL16
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER li1 ;
        RECT 0.590 -13.570 1.010 -13.130 ;
      LAYER mcon ;
        RECT 0.680 -13.480 0.950 -13.210 ;
      LAYER met1 ;
        RECT 0.590 -13.120 1.010 -12.650 ;
        RECT 0.580 -13.570 1.010 -13.120 ;
      LAYER via ;
        RECT 0.680 -12.980 0.950 -12.710 ;
      LAYER met2 ;
        RECT 0.580 -13.120 1.010 -12.610 ;
        RECT 0.590 -13.130 1.010 -13.120 ;
    END
  END WL16
  PIN WL17
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER li1 ;
        RECT 0.590 -14.460 1.010 -14.020 ;
      LAYER mcon ;
        RECT 0.680 -14.380 0.950 -14.110 ;
      LAYER met1 ;
        RECT 0.580 -14.470 1.010 -14.020 ;
        RECT 0.590 -14.940 1.010 -14.470 ;
      LAYER via ;
        RECT 0.680 -14.880 0.950 -14.610 ;
      LAYER met2 ;
        RECT 0.590 -14.980 1.010 -14.450 ;
    END
  END WL17
  PIN WL18
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER li1 ;
        RECT 0.590 -17.180 1.010 -16.740 ;
      LAYER mcon ;
        RECT 0.680 -17.090 0.950 -16.820 ;
      LAYER met1 ;
        RECT 0.590 -16.730 1.010 -16.260 ;
        RECT 0.580 -17.180 1.010 -16.730 ;
      LAYER via ;
        RECT 0.680 -16.590 0.950 -16.320 ;
      LAYER met2 ;
        RECT 0.590 -16.250 1.010 -16.210 ;
        RECT 0.580 -16.730 1.010 -16.250 ;
        RECT 0.590 -16.740 1.010 -16.730 ;
    END
  END WL18
  PIN WL19
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER li1 ;
        RECT 0.590 -18.070 1.010 -17.630 ;
      LAYER mcon ;
        RECT 0.680 -17.990 0.950 -17.720 ;
      LAYER met1 ;
        RECT 0.580 -18.080 1.010 -17.630 ;
        RECT 0.590 -18.550 1.010 -18.080 ;
      LAYER via ;
        RECT 0.680 -18.490 0.950 -18.220 ;
      LAYER met2 ;
        RECT 0.590 -18.090 1.010 -18.060 ;
        RECT 0.580 -18.570 1.010 -18.090 ;
        RECT 0.590 -18.580 1.010 -18.570 ;
    END
  END WL19
  PIN WL20
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER li1 ;
        RECT 0.590 -20.790 1.010 -20.350 ;
      LAYER mcon ;
        RECT 0.680 -20.700 0.950 -20.430 ;
      LAYER met1 ;
        RECT 0.590 -20.340 1.010 -19.870 ;
        RECT 0.580 -20.790 1.010 -20.340 ;
      LAYER via ;
        RECT 0.680 -20.200 0.950 -19.930 ;
      LAYER met2 ;
        RECT 0.580 -20.340 1.010 -19.830 ;
        RECT 0.590 -20.360 1.010 -20.340 ;
    END
  END WL20
  PIN WL21
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER li1 ;
        RECT 0.590 -21.680 1.010 -21.240 ;
      LAYER mcon ;
        RECT 0.680 -21.600 0.950 -21.330 ;
      LAYER met1 ;
        RECT 0.580 -21.690 1.010 -21.240 ;
        RECT 0.590 -22.160 1.010 -21.690 ;
      LAYER via ;
        RECT 0.680 -22.100 0.950 -21.830 ;
      LAYER met2 ;
        RECT 0.590 -21.690 1.010 -21.680 ;
        RECT 0.580 -22.210 1.010 -21.690 ;
    END
  END WL21
  PIN WL22
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER li1 ;
        RECT 0.590 -24.400 1.010 -23.960 ;
      LAYER mcon ;
        RECT 0.680 -24.310 0.950 -24.040 ;
      LAYER met1 ;
        RECT 0.590 -23.950 1.010 -23.480 ;
        RECT 0.580 -24.400 1.010 -23.950 ;
      LAYER via ;
        RECT 0.680 -23.810 0.950 -23.540 ;
      LAYER met2 ;
        RECT 0.590 -23.970 1.010 -23.450 ;
    END
  END WL22
  PIN WL23
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER li1 ;
        RECT 0.590 -25.290 1.010 -24.850 ;
      LAYER mcon ;
        RECT 0.680 -25.210 0.950 -24.940 ;
      LAYER met1 ;
        RECT 0.580 -25.300 1.010 -24.850 ;
        RECT 0.590 -25.770 1.010 -25.300 ;
      LAYER via ;
        RECT 0.680 -25.710 0.950 -25.440 ;
      LAYER met2 ;
        RECT 0.590 -25.310 1.010 -25.290 ;
        RECT 0.580 -25.820 1.010 -25.310 ;
    END
  END WL23
  PIN WL24
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER li1 ;
        RECT 0.590 -28.010 1.010 -27.570 ;
      LAYER mcon ;
        RECT 0.680 -27.920 0.950 -27.650 ;
      LAYER met1 ;
        RECT 0.590 -27.560 1.010 -27.090 ;
        RECT 0.580 -28.010 1.010 -27.560 ;
      LAYER via ;
        RECT 0.680 -27.420 0.950 -27.150 ;
      LAYER met2 ;
        RECT 0.580 -27.550 1.010 -27.040 ;
        RECT 0.590 -27.570 1.010 -27.550 ;
    END
  END WL24
  PIN WL25
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER li1 ;
        RECT 0.590 -28.900 1.010 -28.460 ;
      LAYER mcon ;
        RECT 0.680 -28.820 0.950 -28.550 ;
      LAYER met1 ;
        RECT 0.580 -28.910 1.010 -28.460 ;
        RECT 0.590 -29.380 1.010 -28.910 ;
      LAYER via ;
        RECT 0.680 -29.320 0.950 -29.050 ;
      LAYER met2 ;
        RECT 0.590 -29.410 1.010 -28.890 ;
    END
  END WL25
  PIN WL26
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER li1 ;
        RECT 0.590 -31.620 1.010 -31.180 ;
      LAYER mcon ;
        RECT 0.680 -31.530 0.950 -31.260 ;
      LAYER met1 ;
        RECT 0.590 -31.170 1.010 -30.700 ;
        RECT 0.580 -31.620 1.010 -31.170 ;
      LAYER via ;
        RECT 0.680 -31.030 0.950 -30.760 ;
      LAYER met2 ;
        RECT 0.580 -31.170 1.010 -30.650 ;
        RECT 0.590 -31.180 1.010 -31.170 ;
    END
  END WL26
  PIN WL27
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER li1 ;
        RECT 0.590 -32.510 1.010 -32.070 ;
      LAYER mcon ;
        RECT 0.680 -32.430 0.950 -32.160 ;
      LAYER met1 ;
        RECT 0.580 -32.520 1.010 -32.070 ;
        RECT 0.590 -32.990 1.010 -32.520 ;
      LAYER via ;
        RECT 0.680 -32.930 0.950 -32.660 ;
      LAYER met2 ;
        RECT 0.590 -32.520 1.010 -32.500 ;
        RECT 0.580 -33.030 1.010 -32.520 ;
    END
  END WL27
  PIN WL28
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER li1 ;
        RECT 0.590 -35.230 1.010 -34.790 ;
      LAYER mcon ;
        RECT 0.680 -35.140 0.950 -34.870 ;
      LAYER met1 ;
        RECT 0.590 -34.780 1.010 -34.310 ;
        RECT 0.580 -35.230 1.010 -34.780 ;
      LAYER via ;
        RECT 0.680 -34.640 0.950 -34.370 ;
      LAYER met2 ;
        RECT 0.590 -34.290 1.010 -34.280 ;
        RECT 0.580 -34.770 1.010 -34.290 ;
        RECT 0.590 -34.800 1.010 -34.770 ;
    END
  END WL28
  PIN WL29
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER li1 ;
        RECT 0.590 -36.120 1.010 -35.680 ;
      LAYER mcon ;
        RECT 0.680 -36.040 0.950 -35.770 ;
      LAYER met1 ;
        RECT 0.580 -36.130 1.010 -35.680 ;
        RECT 0.590 -36.600 1.010 -36.130 ;
      LAYER via ;
        RECT 0.680 -36.540 0.950 -36.270 ;
      LAYER met2 ;
        RECT 0.590 -36.130 1.010 -36.120 ;
        RECT 0.580 -36.610 1.010 -36.130 ;
        RECT 0.590 -36.650 1.010 -36.610 ;
    END
  END WL29
  PIN WL30
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER li1 ;
        RECT 0.590 -38.840 1.010 -38.400 ;
      LAYER mcon ;
        RECT 0.680 -38.750 0.950 -38.480 ;
      LAYER met1 ;
        RECT 0.590 -38.390 1.010 -37.920 ;
        RECT 0.580 -38.840 1.010 -38.390 ;
      LAYER via ;
        RECT 0.680 -38.250 0.950 -37.980 ;
      LAYER met2 ;
        RECT 0.590 -38.410 1.010 -37.880 ;
    END
  END WL30
  PIN WL31
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER li1 ;
        RECT 0.590 -39.730 1.010 -39.290 ;
      LAYER mcon ;
        RECT 0.680 -39.650 0.950 -39.380 ;
      LAYER met1 ;
        RECT 0.580 -39.740 1.010 -39.290 ;
        RECT 0.590 -40.210 1.010 -39.740 ;
      LAYER via ;
        RECT 0.680 -40.150 0.950 -39.880 ;
      LAYER met2 ;
        RECT 0.590 -39.740 1.010 -39.730 ;
        RECT 0.580 -40.250 1.010 -39.740 ;
    END
  END WL31
  PIN BL16
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met1 ;
        RECT 109.540 18.860 109.560 18.880 ;
        RECT 109.300 -43.100 109.980 -41.550 ;
    END
  END BL16
  PIN BLb16
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met1 ;
        RECT 114.690 18.780 114.710 18.800 ;
        RECT 114.400 -43.120 115.080 -41.550 ;
    END
  END BLb16
  PIN BL17
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met1 ;
        RECT 116.380 18.740 116.400 18.760 ;
        RECT 116.040 -43.110 116.720 -41.550 ;
    END
  END BL17
  PIN BLb17
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met1 ;
        RECT 121.460 18.750 121.480 18.770 ;
        RECT 121.160 -43.110 121.840 -41.550 ;
    END
  END BLb17
  PIN BL18
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met1 ;
        RECT 123.100 18.790 123.120 18.810 ;
        RECT 122.800 -43.110 123.480 -41.550 ;
    END
  END BL18
  PIN BLb18
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met1 ;
        RECT 128.190 18.710 128.210 18.730 ;
        RECT 127.910 -43.120 128.590 -41.550 ;
    END
  END BLb18
  PIN BL19
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met1 ;
        RECT 129.810 18.630 129.830 18.650 ;
        RECT 129.550 -43.110 130.230 -41.550 ;
    END
  END BL19
  PIN BLb19
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met1 ;
        RECT 134.950 18.810 134.970 18.830 ;
        RECT 134.650 -43.100 135.330 -41.550 ;
    END
  END BLb19
  PIN BL20
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met1 ;
        RECT 136.580 18.730 136.600 18.750 ;
        RECT 136.300 -43.100 136.980 -41.550 ;
    END
  END BL20
  PIN BLb20
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met1 ;
        RECT 141.690 18.750 141.710 18.770 ;
        RECT 141.400 -43.110 142.080 -41.550 ;
    END
  END BLb20
  PIN BL21
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met1 ;
        RECT 143.360 18.700 143.380 18.720 ;
        RECT 143.040 -43.120 143.720 -41.550 ;
    END
  END BL21
  PIN BLb21
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met1 ;
        RECT 148.450 18.780 148.470 18.800 ;
        RECT 148.150 -43.110 148.830 -41.550 ;
    END
  END BLb21
  PIN BL22
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met1 ;
        RECT 150.120 18.760 150.140 18.780 ;
        RECT 149.790 -43.110 150.470 -41.550 ;
    END
  END BL22
  PIN BLb22
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met1 ;
        RECT 155.220 18.720 155.240 18.740 ;
        RECT 154.910 -43.110 155.590 -41.550 ;
    END
  END BLb22
  PIN BL23
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met1 ;
        RECT 156.810 18.770 156.830 18.790 ;
        RECT 156.550 -43.120 157.230 -41.550 ;
    END
  END BL23
  PIN BLb23
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met1 ;
        RECT 162.030 18.780 162.050 18.800 ;
        RECT 161.650 -43.100 162.330 -41.550 ;
    END
  END BLb23
  PIN BL24
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met1 ;
        RECT 163.660 18.730 163.680 18.750 ;
        RECT 163.300 -43.100 163.980 -41.550 ;
    END
  END BL24
  PIN BLb24
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met1 ;
        RECT 168.710 18.640 168.730 18.660 ;
        RECT 168.400 -43.120 169.080 -41.550 ;
    END
  END BLb24
  PIN BL25
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met1 ;
        RECT 170.340 18.650 170.360 18.670 ;
        RECT 170.040 -43.110 170.720 -41.550 ;
    END
  END BL25
  PIN BLb25
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met1 ;
        RECT 175.500 18.800 175.520 18.820 ;
        RECT 175.160 -43.110 175.840 -41.550 ;
    END
  END BLb25
  PIN BL26
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met1 ;
        RECT 177.140 18.690 177.160 18.710 ;
        RECT 176.800 -43.110 177.480 -41.550 ;
    END
  END BL26
  PIN BLb26
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met1 ;
        RECT 182.200 18.670 182.220 18.690 ;
        RECT 181.910 -43.120 182.590 -41.550 ;
    END
  END BLb26
  PIN BL27
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met1 ;
        RECT 183.820 18.780 183.840 18.800 ;
        RECT 183.550 -43.110 184.230 -41.550 ;
    END
  END BL27
  PIN BLb27
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met1 ;
        RECT 188.970 18.790 188.990 18.810 ;
        RECT 188.650 -43.100 189.330 -41.550 ;
    END
  END BLb27
  PIN BL28
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met1 ;
        RECT 190.640 18.750 190.660 18.770 ;
        RECT 190.300 -43.100 190.980 -41.550 ;
    END
  END BL28
  PIN BLb28
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met1 ;
        RECT 195.680 18.730 195.700 18.750 ;
        RECT 195.400 -43.110 196.080 -41.550 ;
    END
  END BLb28
  PIN BL29
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met1 ;
        RECT 197.360 18.810 197.380 18.830 ;
        RECT 197.040 -43.120 197.720 -41.550 ;
    END
  END BL29
  PIN BLb29
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met1 ;
        RECT 202.440 18.680 202.460 18.700 ;
        RECT 202.150 -43.110 202.830 -41.550 ;
    END
  END BLb29
  PIN BL30
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met1 ;
        RECT 204.120 18.710 204.140 18.730 ;
        RECT 203.790 -43.110 204.470 -41.550 ;
    END
  END BL30
  PIN BLb30
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met1 ;
        RECT 209.260 18.700 209.280 18.720 ;
        RECT 208.910 -43.110 209.590 -41.550 ;
    END
  END BLb30
  PIN BL31
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met1 ;
        RECT 210.870 18.710 210.890 18.730 ;
        RECT 210.550 -43.120 211.230 -41.550 ;
    END
  END BL31
  PIN BLb31
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met1 ;
        RECT 215.930 18.650 215.950 18.670 ;
        RECT 215.650 -43.100 216.330 -41.550 ;
    END
  END BLb31
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 3.920 -43.310 4.470 -41.550 ;
        RECT 10.660 -43.350 11.210 -41.550 ;
        RECT 17.420 -43.350 17.970 -41.550 ;
        RECT 24.160 -43.350 24.710 -41.550 ;
        RECT 30.920 -43.350 31.470 -41.550 ;
        RECT 37.660 -43.350 38.210 -41.550 ;
        RECT 44.420 -43.350 44.970 -41.550 ;
        RECT 51.160 -43.310 51.710 -41.550 ;
        RECT 57.920 -43.310 58.470 -41.550 ;
        RECT 64.660 -43.350 65.210 -41.550 ;
        RECT 71.420 -43.350 71.970 -41.550 ;
        RECT 78.160 -43.350 78.710 -41.550 ;
        RECT 84.920 -43.350 85.470 -41.550 ;
        RECT 91.660 -43.350 92.210 -41.550 ;
        RECT 98.420 -43.350 98.970 -41.550 ;
        RECT 105.160 -43.310 105.710 -41.550 ;
        RECT 111.920 -43.310 112.470 -41.550 ;
        RECT 118.660 -43.350 119.210 -41.550 ;
        RECT 125.420 -43.350 125.970 -41.550 ;
        RECT 132.160 -43.350 132.710 -41.550 ;
        RECT 138.920 -43.350 139.470 -41.550 ;
        RECT 145.660 -43.350 146.210 -41.550 ;
        RECT 152.420 -43.350 152.970 -41.550 ;
        RECT 159.160 -43.310 159.710 -41.550 ;
        RECT 165.920 -43.310 166.470 -41.550 ;
        RECT 172.660 -43.350 173.210 -41.550 ;
        RECT 179.420 -43.350 179.970 -41.550 ;
        RECT 186.160 -43.350 186.710 -41.550 ;
        RECT 192.920 -43.350 193.470 -41.550 ;
        RECT 199.660 -43.350 200.210 -41.550 ;
        RECT 206.420 -43.350 206.970 -41.550 ;
        RECT 213.160 -43.310 213.710 -41.550 ;
      LAYER met2 ;
        RECT -0.790 17.920 1.010 18.980 ;
        RECT 219.350 17.920 221.150 18.980 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT -0.050 17.070 1.010 22.400 ;
        RECT -0.060 16.750 1.010 17.070 ;
        RECT 0.600 16.680 1.010 16.750 ;
        RECT 0.600 13.400 1.010 13.500 ;
        RECT 0.390 13.210 1.010 13.400 ;
        RECT 0.600 13.060 1.010 13.210 ;
        RECT 0.600 9.450 1.010 9.890 ;
        RECT 0.600 6.130 1.010 6.280 ;
        RECT 0.390 5.940 1.010 6.130 ;
        RECT 0.600 5.840 1.010 5.940 ;
        RECT 0.600 2.630 1.010 2.670 ;
        RECT -0.060 2.270 1.010 2.630 ;
        RECT 0.600 2.230 1.010 2.270 ;
        RECT 0.600 -1.040 1.010 -0.940 ;
        RECT 0.390 -1.230 1.010 -1.040 ;
        RECT 0.600 -1.380 1.010 -1.230 ;
        RECT 0.600 -4.990 1.010 -4.550 ;
        RECT 0.600 -8.310 1.010 -8.160 ;
        RECT 0.390 -8.500 1.010 -8.310 ;
        RECT 0.600 -8.600 1.010 -8.500 ;
        RECT 0.600 -11.810 1.010 -11.770 ;
        RECT -0.060 -12.170 1.010 -11.810 ;
        RECT 0.600 -12.210 1.010 -12.170 ;
        RECT 0.600 -15.480 1.010 -15.380 ;
        RECT 0.390 -15.670 1.010 -15.480 ;
        RECT 0.600 -15.820 1.010 -15.670 ;
        RECT 0.600 -19.430 1.010 -18.990 ;
        RECT 0.600 -22.750 1.010 -22.600 ;
        RECT 0.390 -22.940 1.010 -22.750 ;
        RECT 0.600 -23.040 1.010 -22.940 ;
        RECT 0.600 -26.250 1.010 -26.210 ;
        RECT -0.060 -26.610 1.010 -26.250 ;
        RECT 0.600 -26.650 1.010 -26.610 ;
        RECT 0.600 -29.920 1.010 -29.820 ;
        RECT 0.390 -30.110 1.010 -29.920 ;
        RECT 0.600 -30.260 1.010 -30.110 ;
        RECT 0.600 -33.870 1.010 -33.430 ;
        RECT 0.600 -37.190 1.010 -37.040 ;
        RECT 0.390 -37.380 1.010 -37.190 ;
        RECT 0.600 -37.480 1.010 -37.380 ;
        RECT 0.600 -40.730 1.010 -40.660 ;
        RECT -0.060 -41.050 1.010 -40.730 ;
        RECT 0.600 -41.090 1.010 -41.050 ;
      LAYER mcon ;
        RECT 0.110 20.190 0.810 22.070 ;
      LAYER met1 ;
        RECT -0.110 22.680 1.150 24.140 ;
        RECT -0.110 22.210 1.010 22.680 ;
        RECT -0.130 20.070 1.010 22.210 ;
        RECT -0.110 20.030 1.010 20.070 ;
      LAYER via ;
        RECT 0.170 22.270 0.830 23.840 ;
      LAYER met2 ;
        RECT -0.680 22.110 1.780 24.480 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 1.010 -41.100 217.690 22.400 ;
      LAYER met1 ;
        RECT 1.010 -41.550 217.050 22.680 ;
      LAYER met2 ;
        RECT 1.010 -40.250 219.350 18.980 ;
  END
END IMPACTSram
END LIBRARY

