VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO IMPACTSram
  CLASS BLOCK ;
  FOREIGN IMPACTSram ;
  ORIGIN 0.790 43.350 ;
  SIZE 221.940 BY 62.720 ;
  PIN BL0
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met1 ;
        RECT 1.660 18.680 1.680 18.700 ;
    END
  END BL0
  PIN BLb0
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met1 ;
        RECT 6.780 18.630 6.800 18.650 ;
    END
  END BLb0
  PIN BL1
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met1 ;
        RECT 8.390 18.590 8.410 18.610 ;
    END
  END BL1
  PIN BLb1
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met1 ;
        RECT 13.540 18.470 13.560 18.490 ;
    END
  END BLb1
  PIN BL2
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met1 ;
        RECT 15.150 18.510 15.170 18.530 ;
    END
  END BL2
  PIN BLb2
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met1 ;
        RECT 20.310 18.700 20.330 18.720 ;
    END
  END BLb2
  PIN BL3
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met1 ;
        RECT 21.870 18.620 21.890 18.640 ;
    END
  END BL3
  PIN BLb3
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met1 ;
        RECT 26.990 18.690 27.010 18.710 ;
    END
  END BLb3
  PIN BL4
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met1 ;
        RECT 28.690 18.720 28.710 18.740 ;
    END
  END BL4
  PIN BLb4
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met1 ;
        RECT 33.780 18.700 33.800 18.720 ;
    END
  END BLb4
  PIN BL5
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met1 ;
        RECT 35.450 18.690 35.470 18.710 ;
    END
  END BL5
  PIN BLb5
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met1 ;
        RECT 40.530 18.460 40.550 18.480 ;
    END
  END BLb5
  PIN BL6
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met1 ;
        RECT 42.170 18.510 42.190 18.530 ;
    END
  END BL6
  PIN BLb6
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met1 ;
        RECT 47.280 18.350 47.300 18.370 ;
    END
  END BLb6
  PIN BL7
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met1 ;
        RECT 48.930 18.780 48.950 18.800 ;
    END
  END BL7
  PIN BLb7
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met1 ;
        RECT 53.970 18.680 53.990 18.700 ;
    END
  END BLb7
  PIN BL8
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met1 ;
        RECT 55.680 18.700 55.700 18.720 ;
    END
  END BL8
  PIN BLb8
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met1 ;
        RECT 60.870 18.720 60.890 18.740 ;
    END
  END BLb8
  PIN BL9
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met1 ;
        RECT 62.410 18.820 62.430 18.840 ;
    END
  END BL9
  PIN BLb9
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met1 ;
        RECT 67.510 18.850 67.530 18.870 ;
    END
  END BLb9
  PIN BL10
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met1 ;
        RECT 69.120 18.820 69.140 18.840 ;
    END
  END BL10
  PIN BLb10
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met1 ;
        RECT 74.310 18.820 74.330 18.840 ;
    END
  END BLb10
  PIN BL11
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met1 ;
        RECT 75.910 18.810 75.930 18.830 ;
    END
  END BL11
  PIN BLb11
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met1 ;
        RECT 81.040 18.890 81.060 18.910 ;
    END
  END BLb11
  PIN BL12
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met1 ;
        RECT 82.640 18.620 82.660 18.640 ;
    END
  END BL12
  PIN BLb12
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met1 ;
        RECT 87.780 18.510 87.800 18.530 ;
    END
  END BLb12
  PIN BL13
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met1 ;
        RECT 89.410 18.560 89.430 18.580 ;
    END
  END BL13
  PIN BLb13
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met1 ;
        RECT 94.530 18.550 94.550 18.570 ;
    END
  END BLb13
  PIN BL14
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met1 ;
        RECT 96.150 18.390 96.170 18.410 ;
    END
  END BL14
  PIN BLb14
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met1 ;
        RECT 101.310 18.490 101.330 18.510 ;
    END
  END BLb14
  PIN BL15
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met1 ;
        RECT 102.870 18.600 102.890 18.620 ;
    END
  END BL15
  PIN BLb15
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met1 ;
        RECT 108.020 18.410 108.040 18.430 ;
    END
  END BLb15
  PIN WL0
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER met2 ;
        RECT 0.740 15.860 0.760 15.880 ;
    END
  END WL0
  PIN WL1
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER met2 ;
        RECT 0.790 14.080 0.810 14.100 ;
    END
  END WL1
  PIN WL2
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER met2 ;
        RECT 0.960 12.230 0.980 12.250 ;
    END
  END WL2
  PIN WL3
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER met2 ;
        RECT 1.040 10.460 1.060 10.480 ;
    END
  END WL3
  PIN WL4
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER met2 ;
        RECT 1.000 8.650 1.020 8.670 ;
    END
  END WL4
  PIN WL5
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER met2 ;
        RECT 1.020 7.100 1.040 7.120 ;
    END
  END WL5
  PIN WL6
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER met2 ;
        RECT 1.050 5.240 1.070 5.260 ;
    END
  END WL6
  PIN WL7
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER met2 ;
        RECT 1.010 3.470 1.030 3.490 ;
    END
  END WL7
  PIN WL8
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER met2 ;
        RECT 1.030 1.590 1.050 1.610 ;
    END
  END WL8
  PIN WL9
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER met2 ;
        RECT 1.050 -0.160 1.070 -0.140 ;
    END
  END WL9
  PIN WL10
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER met2 ;
        RECT 1.030 -1.870 1.050 -1.850 ;
    END
  END WL10
  PIN WL11
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER met2 ;
        RECT 1.020 -3.710 1.040 -3.690 ;
    END
  END WL11
  PIN WL12
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER met2 ;
        RECT 1.010 -5.480 1.030 -5.460 ;
    END
  END WL12
  PIN WL13
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER met2 ;
        RECT 1.030 -7.550 1.050 -7.530 ;
    END
  END WL13
  PIN WL14
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER met2 ;
        RECT 1.010 -9.260 1.030 -9.240 ;
    END
  END WL14
  PIN WL15
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER met2 ;
        RECT 1.010 -10.970 1.030 -10.950 ;
    END
  END WL15
  PIN WL16
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER met2 ;
        RECT 0.930 -12.980 0.950 -12.960 ;
    END
  END WL16
  PIN WL17
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER met2 ;
        RECT 0.930 -14.800 0.950 -14.780 ;
    END
  END WL17
  PIN WL18
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER met2 ;
        RECT 0.830 -16.480 0.850 -16.460 ;
    END
  END WL18
  PIN WL19
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER met2 ;
        RECT 0.850 -18.330 0.870 -18.310 ;
    END
  END WL19
  PIN WL20
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER met2 ;
        RECT 0.790 -20.090 0.810 -20.070 ;
    END
  END WL20
  PIN WL21
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER met2 ;
        RECT 0.780 -22.020 0.800 -22.000 ;
    END
  END WL21
  PIN WL22
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER met2 ;
        RECT 0.780 -23.760 0.800 -23.740 ;
    END
  END WL22
  PIN WL23
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER met2 ;
        RECT 0.810 -25.640 0.830 -25.620 ;
    END
  END WL23
  PIN WL24
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER met2 ;
        RECT 0.790 -27.350 0.810 -27.330 ;
    END
  END WL24
  PIN WL25
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER met2 ;
        RECT 0.800 -29.210 0.820 -29.190 ;
    END
  END WL25
  PIN WL26
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER met2 ;
        RECT 0.800 -30.930 0.820 -30.910 ;
    END
  END WL26
  PIN WL27
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER met2 ;
        RECT 0.790 -32.810 0.810 -32.790 ;
    END
  END WL27
  PIN WL28
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER met2 ;
        RECT 0.790 -34.540 0.810 -34.520 ;
    END
  END WL28
  PIN WL29
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER met2 ;
        RECT 0.800 -36.450 0.820 -36.430 ;
    END
  END WL29
  PIN WL30
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER met2 ;
        RECT 0.780 -38.140 0.800 -38.120 ;
    END
  END WL30
  PIN WL31
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER met2 ;
        RECT 0.790 -40.020 0.810 -40.000 ;
    END
  END WL31
  PIN BL16
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met1 ;
        RECT 109.540 18.860 109.560 18.880 ;
    END
  END BL16
  PIN BLb16
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met1 ;
        RECT 114.690 18.780 114.710 18.800 ;
    END
  END BLb16
  PIN BL17
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met1 ;
        RECT 116.380 18.740 116.400 18.760 ;
    END
  END BL17
  PIN BLb17
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met1 ;
        RECT 121.460 18.750 121.480 18.770 ;
    END
  END BLb17
  PIN BL18
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met1 ;
        RECT 123.100 18.790 123.120 18.810 ;
    END
  END BL18
  PIN BLb18
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met1 ;
        RECT 128.190 18.710 128.210 18.730 ;
    END
  END BLb18
  PIN BL19
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met1 ;
        RECT 129.810 18.630 129.830 18.650 ;
    END
  END BL19
  PIN BLb19
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met1 ;
        RECT 134.950 18.810 134.970 18.830 ;
    END
  END BLb19
  PIN BL20
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met1 ;
        RECT 136.580 18.730 136.600 18.750 ;
    END
  END BL20
  PIN BLb20
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met1 ;
        RECT 141.690 18.750 141.710 18.770 ;
    END
  END BLb20
  PIN BL21
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met1 ;
        RECT 143.360 18.700 143.380 18.720 ;
    END
  END BL21
  PIN BLb21
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met1 ;
        RECT 148.450 18.780 148.470 18.800 ;
    END
  END BLb21
  PIN BL22
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met1 ;
        RECT 150.120 18.760 150.140 18.780 ;
    END
  END BL22
  PIN BLb22
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met1 ;
        RECT 155.220 18.720 155.240 18.740 ;
    END
  END BLb22
  PIN BL23
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met1 ;
        RECT 156.810 18.770 156.830 18.790 ;
    END
  END BL23
  PIN BLb23
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met1 ;
        RECT 162.030 18.780 162.050 18.800 ;
    END
  END BLb23
  PIN BL24
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met1 ;
        RECT 163.660 18.730 163.680 18.750 ;
    END
  END BL24
  PIN BLb24
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met1 ;
        RECT 168.710 18.640 168.730 18.660 ;
    END
  END BLb24
  PIN BL25
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met1 ;
        RECT 170.340 18.650 170.360 18.670 ;
    END
  END BL25
  PIN BLb25
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met1 ;
        RECT 175.500 18.800 175.520 18.820 ;
    END
  END BLb25
  PIN BL26
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met1 ;
        RECT 177.140 18.690 177.160 18.710 ;
    END
  END BL26
  PIN BLb26
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met1 ;
        RECT 182.200 18.670 182.220 18.690 ;
    END
  END BLb26
  PIN BL27
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met1 ;
        RECT 183.820 18.780 183.840 18.800 ;
    END
  END BL27
  PIN BLb27
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met1 ;
        RECT 188.970 18.790 188.990 18.810 ;
    END
  END BLb27
  PIN BL28
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met1 ;
        RECT 190.640 18.750 190.660 18.770 ;
    END
  END BL28
  PIN BLb28
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met1 ;
        RECT 195.680 18.730 195.700 18.750 ;
    END
  END BLb28
  PIN BL29
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met1 ;
        RECT 197.360 18.810 197.380 18.830 ;
    END
  END BL29
  PIN BLb29
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met1 ;
        RECT 202.440 18.680 202.460 18.700 ;
    END
  END BLb29
  PIN BL30
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met1 ;
        RECT 204.120 18.710 204.140 18.730 ;
    END
  END BL30
  PIN BLb30
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met1 ;
        RECT 209.260 18.700 209.280 18.720 ;
    END
  END BLb30
  PIN BL31
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met1 ;
        RECT 210.870 18.710 210.890 18.730 ;
    END
  END BL31
  PIN BLb31
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met1 ;
        RECT 215.930 18.650 215.950 18.670 ;
    END
  END BLb31
  PIN VPWR
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 0.120 18.430 0.130 18.440 ;
    END
  END VPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.300 16.900 0.310 16.910 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT -0.060 17.080 217.690 17.120 ;
        RECT -0.060 16.730 0.130 17.080 ;
        RECT 0.480 16.730 217.690 17.080 ;
        RECT -0.060 -41.100 217.690 16.730 ;
      LAYER met1 ;
        RECT 0.580 19.190 217.050 19.370 ;
        RECT 0.580 19.150 80.760 19.190 ;
        RECT 0.580 19.120 67.230 19.150 ;
        RECT 0.580 19.080 62.130 19.120 ;
        RECT 0.580 19.020 48.650 19.080 ;
        RECT 0.580 19.000 28.410 19.020 ;
        RECT 0.580 18.980 20.030 19.000 ;
        RECT 0.580 18.400 1.380 18.980 ;
        RECT 1.960 18.930 20.030 18.980 ;
        RECT 1.960 18.400 6.500 18.930 ;
        RECT 0.580 18.350 6.500 18.400 ;
        RECT 7.080 18.890 20.030 18.930 ;
        RECT 7.080 18.350 8.110 18.890 ;
        RECT 0.580 18.310 8.110 18.350 ;
        RECT 8.690 18.810 20.030 18.890 ;
        RECT 8.690 18.770 14.870 18.810 ;
        RECT 8.690 18.310 13.260 18.770 ;
        RECT 0.580 18.190 13.260 18.310 ;
        RECT 13.840 18.230 14.870 18.770 ;
        RECT 15.450 18.420 20.030 18.810 ;
        RECT 20.610 18.990 28.410 19.000 ;
        RECT 20.610 18.920 26.710 18.990 ;
        RECT 20.610 18.420 21.590 18.920 ;
        RECT 15.450 18.340 21.590 18.420 ;
        RECT 22.170 18.410 26.710 18.920 ;
        RECT 27.290 18.440 28.410 18.990 ;
        RECT 28.990 19.000 48.650 19.020 ;
        RECT 28.990 18.440 33.500 19.000 ;
        RECT 27.290 18.420 33.500 18.440 ;
        RECT 34.080 18.990 48.650 19.000 ;
        RECT 34.080 18.420 35.170 18.990 ;
        RECT 27.290 18.410 35.170 18.420 ;
        RECT 35.750 18.810 48.650 18.990 ;
        RECT 35.750 18.760 41.890 18.810 ;
        RECT 35.750 18.410 40.250 18.760 ;
        RECT 22.170 18.340 40.250 18.410 ;
        RECT 15.450 18.230 40.250 18.340 ;
        RECT 13.840 18.190 40.250 18.230 ;
        RECT 0.580 18.180 40.250 18.190 ;
        RECT 40.830 18.230 41.890 18.760 ;
        RECT 42.470 18.650 48.650 18.810 ;
        RECT 42.470 18.230 47.000 18.650 ;
        RECT 40.830 18.180 47.000 18.230 ;
        RECT 0.580 18.070 47.000 18.180 ;
        RECT 47.580 18.500 48.650 18.650 ;
        RECT 49.230 19.020 62.130 19.080 ;
        RECT 49.230 19.000 60.590 19.020 ;
        RECT 49.230 18.980 55.400 19.000 ;
        RECT 49.230 18.500 53.690 18.980 ;
        RECT 47.580 18.400 53.690 18.500 ;
        RECT 54.270 18.420 55.400 18.980 ;
        RECT 55.980 18.440 60.590 19.000 ;
        RECT 61.170 18.540 62.130 19.020 ;
        RECT 62.710 18.570 67.230 19.120 ;
        RECT 67.810 19.120 80.760 19.150 ;
        RECT 67.810 18.570 68.840 19.120 ;
        RECT 62.710 18.540 68.840 18.570 ;
        RECT 69.420 18.540 74.030 19.120 ;
        RECT 74.610 19.110 80.760 19.120 ;
        RECT 74.610 18.540 75.630 19.110 ;
        RECT 61.170 18.530 75.630 18.540 ;
        RECT 76.210 18.610 80.760 19.110 ;
        RECT 81.340 19.160 217.050 19.190 ;
        RECT 81.340 18.920 109.260 19.160 ;
        RECT 81.340 18.610 82.360 18.920 ;
        RECT 76.210 18.530 82.360 18.610 ;
        RECT 61.170 18.440 82.360 18.530 ;
        RECT 55.980 18.420 82.360 18.440 ;
        RECT 54.270 18.400 82.360 18.420 ;
        RECT 47.580 18.340 82.360 18.400 ;
        RECT 82.940 18.900 109.260 18.920 ;
        RECT 82.940 18.860 102.590 18.900 ;
        RECT 82.940 18.810 89.130 18.860 ;
        RECT 82.940 18.340 87.500 18.810 ;
        RECT 47.580 18.230 87.500 18.340 ;
        RECT 88.080 18.280 89.130 18.810 ;
        RECT 89.710 18.850 102.590 18.860 ;
        RECT 89.710 18.280 94.250 18.850 ;
        RECT 88.080 18.270 94.250 18.280 ;
        RECT 94.830 18.790 102.590 18.850 ;
        RECT 94.830 18.690 101.030 18.790 ;
        RECT 94.830 18.270 95.870 18.690 ;
        RECT 88.080 18.230 95.870 18.270 ;
        RECT 47.580 18.110 95.870 18.230 ;
        RECT 96.450 18.210 101.030 18.690 ;
        RECT 101.610 18.320 102.590 18.790 ;
        RECT 103.170 18.710 109.260 18.900 ;
        RECT 103.170 18.320 107.740 18.710 ;
        RECT 101.610 18.210 107.740 18.320 ;
        RECT 96.450 18.130 107.740 18.210 ;
        RECT 108.320 18.580 109.260 18.710 ;
        RECT 109.840 19.110 217.050 19.160 ;
        RECT 109.840 19.090 134.670 19.110 ;
        RECT 109.840 19.080 122.820 19.090 ;
        RECT 109.840 18.580 114.410 19.080 ;
        RECT 108.320 18.500 114.410 18.580 ;
        RECT 114.990 19.050 122.820 19.080 ;
        RECT 114.990 19.040 121.180 19.050 ;
        RECT 114.990 18.500 116.100 19.040 ;
        RECT 108.320 18.460 116.100 18.500 ;
        RECT 116.680 18.470 121.180 19.040 ;
        RECT 121.760 18.510 122.820 19.050 ;
        RECT 123.400 19.010 134.670 19.090 ;
        RECT 123.400 18.510 127.910 19.010 ;
        RECT 121.760 18.470 127.910 18.510 ;
        RECT 116.680 18.460 127.910 18.470 ;
        RECT 108.320 18.430 127.910 18.460 ;
        RECT 128.490 18.930 134.670 19.010 ;
        RECT 128.490 18.430 129.530 18.930 ;
        RECT 108.320 18.350 129.530 18.430 ;
        RECT 130.110 18.530 134.670 18.930 ;
        RECT 135.250 19.100 197.080 19.110 ;
        RECT 135.250 19.080 175.220 19.100 ;
        RECT 135.250 19.050 148.170 19.080 ;
        RECT 135.250 19.030 141.410 19.050 ;
        RECT 135.250 18.530 136.300 19.030 ;
        RECT 130.110 18.450 136.300 18.530 ;
        RECT 136.880 18.470 141.410 19.030 ;
        RECT 141.990 19.000 148.170 19.050 ;
        RECT 141.990 18.470 143.080 19.000 ;
        RECT 136.880 18.450 143.080 18.470 ;
        RECT 130.110 18.420 143.080 18.450 ;
        RECT 143.660 18.500 148.170 19.000 ;
        RECT 148.750 19.070 161.750 19.080 ;
        RECT 148.750 19.060 156.530 19.070 ;
        RECT 148.750 18.500 149.840 19.060 ;
        RECT 143.660 18.480 149.840 18.500 ;
        RECT 150.420 19.020 156.530 19.060 ;
        RECT 150.420 18.480 154.940 19.020 ;
        RECT 143.660 18.440 154.940 18.480 ;
        RECT 155.520 18.490 156.530 19.020 ;
        RECT 157.110 18.500 161.750 19.070 ;
        RECT 162.330 19.030 175.220 19.080 ;
        RECT 162.330 18.500 163.380 19.030 ;
        RECT 157.110 18.490 163.380 18.500 ;
        RECT 155.520 18.450 163.380 18.490 ;
        RECT 163.960 18.950 175.220 19.030 ;
        RECT 163.960 18.940 170.060 18.950 ;
        RECT 163.960 18.450 168.430 18.940 ;
        RECT 155.520 18.440 168.430 18.450 ;
        RECT 143.660 18.420 168.430 18.440 ;
        RECT 130.110 18.360 168.430 18.420 ;
        RECT 169.010 18.370 170.060 18.940 ;
        RECT 170.640 18.520 175.220 18.950 ;
        RECT 175.800 19.090 197.080 19.100 ;
        RECT 175.800 19.080 188.690 19.090 ;
        RECT 175.800 18.990 183.540 19.080 ;
        RECT 175.800 18.520 176.860 18.990 ;
        RECT 170.640 18.410 176.860 18.520 ;
        RECT 177.440 18.970 183.540 18.990 ;
        RECT 177.440 18.410 181.920 18.970 ;
        RECT 170.640 18.390 181.920 18.410 ;
        RECT 182.500 18.500 183.540 18.970 ;
        RECT 184.120 18.510 188.690 19.080 ;
        RECT 189.270 19.050 197.080 19.090 ;
        RECT 189.270 18.510 190.360 19.050 ;
        RECT 184.120 18.500 190.360 18.510 ;
        RECT 182.500 18.470 190.360 18.500 ;
        RECT 190.940 19.030 197.080 19.050 ;
        RECT 190.940 18.470 195.400 19.030 ;
        RECT 182.500 18.450 195.400 18.470 ;
        RECT 195.980 18.530 197.080 19.030 ;
        RECT 197.660 19.010 217.050 19.110 ;
        RECT 197.660 18.980 203.840 19.010 ;
        RECT 197.660 18.530 202.160 18.980 ;
        RECT 195.980 18.450 202.160 18.530 ;
        RECT 182.500 18.400 202.160 18.450 ;
        RECT 202.740 18.430 203.840 18.980 ;
        RECT 204.420 19.000 210.590 19.010 ;
        RECT 204.420 18.430 208.980 19.000 ;
        RECT 202.740 18.420 208.980 18.430 ;
        RECT 209.560 18.430 210.590 19.000 ;
        RECT 211.170 18.950 217.050 19.010 ;
        RECT 211.170 18.430 215.650 18.950 ;
        RECT 209.560 18.420 215.650 18.430 ;
        RECT 202.740 18.400 215.650 18.420 ;
        RECT 182.500 18.390 215.650 18.400 ;
        RECT 170.640 18.370 215.650 18.390 ;
        RECT 216.230 18.370 217.050 18.950 ;
        RECT 169.010 18.360 217.050 18.370 ;
        RECT 130.110 18.350 217.050 18.360 ;
        RECT 108.320 18.130 217.050 18.350 ;
        RECT 96.450 18.110 217.050 18.130 ;
        RECT 47.580 18.070 217.050 18.110 ;
        RECT 0.580 -43.350 217.050 18.070 ;
      LAYER met2 ;
        RECT -0.790 18.440 221.150 18.980 ;
        RECT -0.790 18.430 0.120 18.440 ;
        RECT 0.410 18.430 221.150 18.440 ;
        RECT -0.790 16.160 221.150 18.430 ;
        RECT -0.790 15.580 0.460 16.160 ;
        RECT 1.040 15.580 221.150 16.160 ;
        RECT -0.790 14.380 221.150 15.580 ;
        RECT -0.790 13.800 0.510 14.380 ;
        RECT 1.090 13.800 221.150 14.380 ;
        RECT -0.790 12.530 221.150 13.800 ;
        RECT -0.790 11.950 0.680 12.530 ;
        RECT 1.260 11.950 221.150 12.530 ;
        RECT -0.790 10.760 221.150 11.950 ;
        RECT -0.790 10.180 0.760 10.760 ;
        RECT 1.340 10.180 221.150 10.760 ;
        RECT -0.790 8.950 221.150 10.180 ;
        RECT -0.790 8.370 0.720 8.950 ;
        RECT 1.300 8.370 221.150 8.950 ;
        RECT -0.790 7.400 221.150 8.370 ;
        RECT -0.790 6.820 0.740 7.400 ;
        RECT 1.320 6.820 221.150 7.400 ;
        RECT -0.790 5.540 221.150 6.820 ;
        RECT -0.790 4.960 0.770 5.540 ;
        RECT 1.350 4.960 221.150 5.540 ;
        RECT -0.790 3.770 221.150 4.960 ;
        RECT -0.790 3.190 0.730 3.770 ;
        RECT 1.310 3.190 221.150 3.770 ;
        RECT -0.790 1.890 221.150 3.190 ;
        RECT -0.790 1.310 0.750 1.890 ;
        RECT 1.330 1.310 221.150 1.890 ;
        RECT -0.790 0.140 221.150 1.310 ;
        RECT -0.790 -0.440 0.770 0.140 ;
        RECT 1.350 -0.440 221.150 0.140 ;
        RECT -0.790 -1.570 221.150 -0.440 ;
        RECT -0.790 -2.150 0.750 -1.570 ;
        RECT 1.330 -2.150 221.150 -1.570 ;
        RECT -0.790 -3.410 221.150 -2.150 ;
        RECT -0.790 -3.990 0.740 -3.410 ;
        RECT 1.320 -3.990 221.150 -3.410 ;
        RECT -0.790 -5.180 221.150 -3.990 ;
        RECT -0.790 -5.760 0.730 -5.180 ;
        RECT 1.310 -5.760 221.150 -5.180 ;
        RECT -0.790 -7.250 221.150 -5.760 ;
        RECT -0.790 -7.830 0.750 -7.250 ;
        RECT 1.330 -7.830 221.150 -7.250 ;
        RECT -0.790 -8.960 221.150 -7.830 ;
        RECT -0.790 -9.540 0.730 -8.960 ;
        RECT 1.310 -9.540 221.150 -8.960 ;
        RECT -0.790 -10.670 221.150 -9.540 ;
        RECT -0.790 -11.250 0.730 -10.670 ;
        RECT 1.310 -11.250 221.150 -10.670 ;
        RECT -0.790 -12.680 221.150 -11.250 ;
        RECT -0.790 -13.260 0.650 -12.680 ;
        RECT 1.230 -13.260 221.150 -12.680 ;
        RECT -0.790 -14.500 221.150 -13.260 ;
        RECT -0.790 -15.080 0.650 -14.500 ;
        RECT 1.230 -15.080 221.150 -14.500 ;
        RECT -0.790 -16.180 221.150 -15.080 ;
        RECT -0.790 -16.760 0.550 -16.180 ;
        RECT 1.130 -16.760 221.150 -16.180 ;
        RECT -0.790 -18.030 221.150 -16.760 ;
        RECT -0.790 -18.610 0.570 -18.030 ;
        RECT 1.150 -18.610 221.150 -18.030 ;
        RECT -0.790 -19.790 221.150 -18.610 ;
        RECT -0.790 -20.370 0.510 -19.790 ;
        RECT 1.090 -20.370 221.150 -19.790 ;
        RECT -0.790 -21.720 221.150 -20.370 ;
        RECT -0.790 -22.300 0.500 -21.720 ;
        RECT 1.080 -22.300 221.150 -21.720 ;
        RECT -0.790 -23.460 221.150 -22.300 ;
        RECT -0.790 -24.040 0.500 -23.460 ;
        RECT 1.080 -24.040 221.150 -23.460 ;
        RECT -0.790 -25.340 221.150 -24.040 ;
        RECT -0.790 -25.920 0.530 -25.340 ;
        RECT 1.110 -25.920 221.150 -25.340 ;
        RECT -0.790 -27.050 221.150 -25.920 ;
        RECT -0.790 -27.630 0.510 -27.050 ;
        RECT 1.090 -27.630 221.150 -27.050 ;
        RECT -0.790 -28.910 221.150 -27.630 ;
        RECT -0.790 -29.490 0.520 -28.910 ;
        RECT 1.100 -29.490 221.150 -28.910 ;
        RECT -0.790 -30.630 221.150 -29.490 ;
        RECT -0.790 -31.210 0.520 -30.630 ;
        RECT 1.100 -31.210 221.150 -30.630 ;
        RECT -0.790 -32.510 221.150 -31.210 ;
        RECT -0.790 -33.090 0.510 -32.510 ;
        RECT 1.090 -33.090 221.150 -32.510 ;
        RECT -0.790 -34.240 221.150 -33.090 ;
        RECT -0.790 -34.820 0.510 -34.240 ;
        RECT 1.090 -34.820 221.150 -34.240 ;
        RECT -0.790 -36.150 221.150 -34.820 ;
        RECT -0.790 -36.730 0.520 -36.150 ;
        RECT 1.100 -36.730 221.150 -36.150 ;
        RECT -0.790 -37.840 221.150 -36.730 ;
        RECT -0.790 -38.420 0.500 -37.840 ;
        RECT 1.080 -38.420 221.150 -37.840 ;
        RECT -0.790 -39.720 221.150 -38.420 ;
        RECT -0.790 -40.250 0.510 -39.720 ;
        RECT 1.090 -40.250 221.150 -39.720 ;
  END
END IMPACTSram
END LIBRARY

