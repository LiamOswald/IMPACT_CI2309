VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO IMPACTSram
  CLASS BLOCK ;
  FOREIGN IMPACTSram ;
  ORIGIN 0.000 0.000 ;
  SIZE 800.000 BY 2400.000 ;
  PIN Address[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 156.440 800.000 157.040 ;
    END
  END Address[0]
  PIN Address[1000]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2147.480 4.000 2148.080 ;
    END
  END Address[1000]
  PIN Address[1001]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2151.560 4.000 2152.160 ;
    END
  END Address[1001]
  PIN Address[1002]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2155.640 4.000 2156.240 ;
    END
  END Address[1002]
  PIN Address[1003]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2159.720 4.000 2160.320 ;
    END
  END Address[1003]
  PIN Address[1004]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2163.800 4.000 2164.400 ;
    END
  END Address[1004]
  PIN Address[1005]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2167.880 4.000 2168.480 ;
    END
  END Address[1005]
  PIN Address[1006]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2171.960 4.000 2172.560 ;
    END
  END Address[1006]
  PIN Address[1007]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2176.040 4.000 2176.640 ;
    END
  END Address[1007]
  PIN Address[1008]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2180.120 4.000 2180.720 ;
    END
  END Address[1008]
  PIN Address[1009]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2184.200 4.000 2184.800 ;
    END
  END Address[1009]
  PIN Address[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 564.440 800.000 565.040 ;
    END
  END Address[100]
  PIN Address[1010]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2188.280 4.000 2188.880 ;
    END
  END Address[1010]
  PIN Address[1011]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2192.360 4.000 2192.960 ;
    END
  END Address[1011]
  PIN Address[1012]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2196.440 4.000 2197.040 ;
    END
  END Address[1012]
  PIN Address[1013]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2200.520 4.000 2201.120 ;
    END
  END Address[1013]
  PIN Address[1014]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2204.600 4.000 2205.200 ;
    END
  END Address[1014]
  PIN Address[1015]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2208.680 4.000 2209.280 ;
    END
  END Address[1015]
  PIN Address[1016]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2212.760 4.000 2213.360 ;
    END
  END Address[1016]
  PIN Address[1017]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2216.840 4.000 2217.440 ;
    END
  END Address[1017]
  PIN Address[1018]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2220.920 4.000 2221.520 ;
    END
  END Address[1018]
  PIN Address[1019]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2225.000 4.000 2225.600 ;
    END
  END Address[1019]
  PIN Address[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 568.520 800.000 569.120 ;
    END
  END Address[101]
  PIN Address[1020]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2229.080 4.000 2229.680 ;
    END
  END Address[1020]
  PIN Address[1021]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2233.160 4.000 2233.760 ;
    END
  END Address[1021]
  PIN Address[1022]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2237.240 4.000 2237.840 ;
    END
  END Address[1022]
  PIN Address[1023]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2241.320 4.000 2241.920 ;
    END
  END Address[1023]
  PIN Address[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 572.600 800.000 573.200 ;
    END
  END Address[102]
  PIN Address[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 576.680 800.000 577.280 ;
    END
  END Address[103]
  PIN Address[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 580.760 800.000 581.360 ;
    END
  END Address[104]
  PIN Address[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 584.840 800.000 585.440 ;
    END
  END Address[105]
  PIN Address[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 588.920 800.000 589.520 ;
    END
  END Address[106]
  PIN Address[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 593.000 800.000 593.600 ;
    END
  END Address[107]
  PIN Address[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 597.080 800.000 597.680 ;
    END
  END Address[108]
  PIN Address[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 601.160 800.000 601.760 ;
    END
  END Address[109]
  PIN Address[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 197.240 800.000 197.840 ;
    END
  END Address[10]
  PIN Address[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 605.240 800.000 605.840 ;
    END
  END Address[110]
  PIN Address[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 609.320 800.000 609.920 ;
    END
  END Address[111]
  PIN Address[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 613.400 800.000 614.000 ;
    END
  END Address[112]
  PIN Address[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 617.480 800.000 618.080 ;
    END
  END Address[113]
  PIN Address[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 621.560 800.000 622.160 ;
    END
  END Address[114]
  PIN Address[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 625.640 800.000 626.240 ;
    END
  END Address[115]
  PIN Address[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 629.720 800.000 630.320 ;
    END
  END Address[116]
  PIN Address[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 633.800 800.000 634.400 ;
    END
  END Address[117]
  PIN Address[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 637.880 800.000 638.480 ;
    END
  END Address[118]
  PIN Address[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 641.960 800.000 642.560 ;
    END
  END Address[119]
  PIN Address[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 201.320 800.000 201.920 ;
    END
  END Address[11]
  PIN Address[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 646.040 800.000 646.640 ;
    END
  END Address[120]
  PIN Address[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 650.120 800.000 650.720 ;
    END
  END Address[121]
  PIN Address[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 654.200 800.000 654.800 ;
    END
  END Address[122]
  PIN Address[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 658.280 800.000 658.880 ;
    END
  END Address[123]
  PIN Address[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 662.360 800.000 662.960 ;
    END
  END Address[124]
  PIN Address[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 666.440 800.000 667.040 ;
    END
  END Address[125]
  PIN Address[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 670.520 800.000 671.120 ;
    END
  END Address[126]
  PIN Address[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 674.600 800.000 675.200 ;
    END
  END Address[127]
  PIN Address[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 678.680 800.000 679.280 ;
    END
  END Address[128]
  PIN Address[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 682.760 800.000 683.360 ;
    END
  END Address[129]
  PIN Address[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 205.400 800.000 206.000 ;
    END
  END Address[12]
  PIN Address[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 686.840 800.000 687.440 ;
    END
  END Address[130]
  PIN Address[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 690.920 800.000 691.520 ;
    END
  END Address[131]
  PIN Address[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 695.000 800.000 695.600 ;
    END
  END Address[132]
  PIN Address[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 699.080 800.000 699.680 ;
    END
  END Address[133]
  PIN Address[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 703.160 800.000 703.760 ;
    END
  END Address[134]
  PIN Address[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 707.240 800.000 707.840 ;
    END
  END Address[135]
  PIN Address[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 711.320 800.000 711.920 ;
    END
  END Address[136]
  PIN Address[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 715.400 800.000 716.000 ;
    END
  END Address[137]
  PIN Address[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 719.480 800.000 720.080 ;
    END
  END Address[138]
  PIN Address[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 723.560 800.000 724.160 ;
    END
  END Address[139]
  PIN Address[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 209.480 800.000 210.080 ;
    END
  END Address[13]
  PIN Address[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 727.640 800.000 728.240 ;
    END
  END Address[140]
  PIN Address[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 731.720 800.000 732.320 ;
    END
  END Address[141]
  PIN Address[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 735.800 800.000 736.400 ;
    END
  END Address[142]
  PIN Address[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 739.880 800.000 740.480 ;
    END
  END Address[143]
  PIN Address[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 743.960 800.000 744.560 ;
    END
  END Address[144]
  PIN Address[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 748.040 800.000 748.640 ;
    END
  END Address[145]
  PIN Address[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 752.120 800.000 752.720 ;
    END
  END Address[146]
  PIN Address[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 756.200 800.000 756.800 ;
    END
  END Address[147]
  PIN Address[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 760.280 800.000 760.880 ;
    END
  END Address[148]
  PIN Address[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 764.360 800.000 764.960 ;
    END
  END Address[149]
  PIN Address[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 213.560 800.000 214.160 ;
    END
  END Address[14]
  PIN Address[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 768.440 800.000 769.040 ;
    END
  END Address[150]
  PIN Address[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 772.520 800.000 773.120 ;
    END
  END Address[151]
  PIN Address[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 776.600 800.000 777.200 ;
    END
  END Address[152]
  PIN Address[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 780.680 800.000 781.280 ;
    END
  END Address[153]
  PIN Address[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 784.760 800.000 785.360 ;
    END
  END Address[154]
  PIN Address[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 788.840 800.000 789.440 ;
    END
  END Address[155]
  PIN Address[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 792.920 800.000 793.520 ;
    END
  END Address[156]
  PIN Address[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 797.000 800.000 797.600 ;
    END
  END Address[157]
  PIN Address[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 801.080 800.000 801.680 ;
    END
  END Address[158]
  PIN Address[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 805.160 800.000 805.760 ;
    END
  END Address[159]
  PIN Address[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 217.640 800.000 218.240 ;
    END
  END Address[15]
  PIN Address[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 809.240 800.000 809.840 ;
    END
  END Address[160]
  PIN Address[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 813.320 800.000 813.920 ;
    END
  END Address[161]
  PIN Address[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 817.400 800.000 818.000 ;
    END
  END Address[162]
  PIN Address[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 821.480 800.000 822.080 ;
    END
  END Address[163]
  PIN Address[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 825.560 800.000 826.160 ;
    END
  END Address[164]
  PIN Address[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 829.640 800.000 830.240 ;
    END
  END Address[165]
  PIN Address[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 833.720 800.000 834.320 ;
    END
  END Address[166]
  PIN Address[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 837.800 800.000 838.400 ;
    END
  END Address[167]
  PIN Address[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 841.880 800.000 842.480 ;
    END
  END Address[168]
  PIN Address[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 845.960 800.000 846.560 ;
    END
  END Address[169]
  PIN Address[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 221.720 800.000 222.320 ;
    END
  END Address[16]
  PIN Address[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 850.040 800.000 850.640 ;
    END
  END Address[170]
  PIN Address[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 854.120 800.000 854.720 ;
    END
  END Address[171]
  PIN Address[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 858.200 800.000 858.800 ;
    END
  END Address[172]
  PIN Address[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 862.280 800.000 862.880 ;
    END
  END Address[173]
  PIN Address[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 866.360 800.000 866.960 ;
    END
  END Address[174]
  PIN Address[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 870.440 800.000 871.040 ;
    END
  END Address[175]
  PIN Address[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 874.520 800.000 875.120 ;
    END
  END Address[176]
  PIN Address[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 878.600 800.000 879.200 ;
    END
  END Address[177]
  PIN Address[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 882.680 800.000 883.280 ;
    END
  END Address[178]
  PIN Address[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 886.760 800.000 887.360 ;
    END
  END Address[179]
  PIN Address[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 225.800 800.000 226.400 ;
    END
  END Address[17]
  PIN Address[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 890.840 800.000 891.440 ;
    END
  END Address[180]
  PIN Address[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 894.920 800.000 895.520 ;
    END
  END Address[181]
  PIN Address[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 899.000 800.000 899.600 ;
    END
  END Address[182]
  PIN Address[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 903.080 800.000 903.680 ;
    END
  END Address[183]
  PIN Address[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 907.160 800.000 907.760 ;
    END
  END Address[184]
  PIN Address[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 911.240 800.000 911.840 ;
    END
  END Address[185]
  PIN Address[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 915.320 800.000 915.920 ;
    END
  END Address[186]
  PIN Address[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 919.400 800.000 920.000 ;
    END
  END Address[187]
  PIN Address[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 923.480 800.000 924.080 ;
    END
  END Address[188]
  PIN Address[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 927.560 800.000 928.160 ;
    END
  END Address[189]
  PIN Address[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 229.880 800.000 230.480 ;
    END
  END Address[18]
  PIN Address[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 931.640 800.000 932.240 ;
    END
  END Address[190]
  PIN Address[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 935.720 800.000 936.320 ;
    END
  END Address[191]
  PIN Address[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 939.800 800.000 940.400 ;
    END
  END Address[192]
  PIN Address[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 943.880 800.000 944.480 ;
    END
  END Address[193]
  PIN Address[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 947.960 800.000 948.560 ;
    END
  END Address[194]
  PIN Address[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 952.040 800.000 952.640 ;
    END
  END Address[195]
  PIN Address[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 956.120 800.000 956.720 ;
    END
  END Address[196]
  PIN Address[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 960.200 800.000 960.800 ;
    END
  END Address[197]
  PIN Address[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 964.280 800.000 964.880 ;
    END
  END Address[198]
  PIN Address[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 968.360 800.000 968.960 ;
    END
  END Address[199]
  PIN Address[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 233.960 800.000 234.560 ;
    END
  END Address[19]
  PIN Address[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 160.520 800.000 161.120 ;
    END
  END Address[1]
  PIN Address[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 972.440 800.000 973.040 ;
    END
  END Address[200]
  PIN Address[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 976.520 800.000 977.120 ;
    END
  END Address[201]
  PIN Address[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 980.600 800.000 981.200 ;
    END
  END Address[202]
  PIN Address[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 984.680 800.000 985.280 ;
    END
  END Address[203]
  PIN Address[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 988.760 800.000 989.360 ;
    END
  END Address[204]
  PIN Address[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 992.840 800.000 993.440 ;
    END
  END Address[205]
  PIN Address[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 996.920 800.000 997.520 ;
    END
  END Address[206]
  PIN Address[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1001.000 800.000 1001.600 ;
    END
  END Address[207]
  PIN Address[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1005.080 800.000 1005.680 ;
    END
  END Address[208]
  PIN Address[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1009.160 800.000 1009.760 ;
    END
  END Address[209]
  PIN Address[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 238.040 800.000 238.640 ;
    END
  END Address[20]
  PIN Address[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1013.240 800.000 1013.840 ;
    END
  END Address[210]
  PIN Address[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1017.320 800.000 1017.920 ;
    END
  END Address[211]
  PIN Address[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1021.400 800.000 1022.000 ;
    END
  END Address[212]
  PIN Address[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1025.480 800.000 1026.080 ;
    END
  END Address[213]
  PIN Address[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1029.560 800.000 1030.160 ;
    END
  END Address[214]
  PIN Address[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1033.640 800.000 1034.240 ;
    END
  END Address[215]
  PIN Address[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1037.720 800.000 1038.320 ;
    END
  END Address[216]
  PIN Address[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1041.800 800.000 1042.400 ;
    END
  END Address[217]
  PIN Address[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1045.880 800.000 1046.480 ;
    END
  END Address[218]
  PIN Address[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1049.960 800.000 1050.560 ;
    END
  END Address[219]
  PIN Address[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 242.120 800.000 242.720 ;
    END
  END Address[21]
  PIN Address[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1054.040 800.000 1054.640 ;
    END
  END Address[220]
  PIN Address[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1058.120 800.000 1058.720 ;
    END
  END Address[221]
  PIN Address[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1062.200 800.000 1062.800 ;
    END
  END Address[222]
  PIN Address[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1066.280 800.000 1066.880 ;
    END
  END Address[223]
  PIN Address[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1070.360 800.000 1070.960 ;
    END
  END Address[224]
  PIN Address[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1074.440 800.000 1075.040 ;
    END
  END Address[225]
  PIN Address[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1078.520 800.000 1079.120 ;
    END
  END Address[226]
  PIN Address[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1082.600 800.000 1083.200 ;
    END
  END Address[227]
  PIN Address[228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1086.680 800.000 1087.280 ;
    END
  END Address[228]
  PIN Address[229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1090.760 800.000 1091.360 ;
    END
  END Address[229]
  PIN Address[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 246.200 800.000 246.800 ;
    END
  END Address[22]
  PIN Address[230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1094.840 800.000 1095.440 ;
    END
  END Address[230]
  PIN Address[231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1098.920 800.000 1099.520 ;
    END
  END Address[231]
  PIN Address[232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1103.000 800.000 1103.600 ;
    END
  END Address[232]
  PIN Address[233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1107.080 800.000 1107.680 ;
    END
  END Address[233]
  PIN Address[234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1111.160 800.000 1111.760 ;
    END
  END Address[234]
  PIN Address[235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1115.240 800.000 1115.840 ;
    END
  END Address[235]
  PIN Address[236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1119.320 800.000 1119.920 ;
    END
  END Address[236]
  PIN Address[237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1123.400 800.000 1124.000 ;
    END
  END Address[237]
  PIN Address[238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1127.480 800.000 1128.080 ;
    END
  END Address[238]
  PIN Address[239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1131.560 800.000 1132.160 ;
    END
  END Address[239]
  PIN Address[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 250.280 800.000 250.880 ;
    END
  END Address[23]
  PIN Address[240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1135.640 800.000 1136.240 ;
    END
  END Address[240]
  PIN Address[241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1139.720 800.000 1140.320 ;
    END
  END Address[241]
  PIN Address[242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1143.800 800.000 1144.400 ;
    END
  END Address[242]
  PIN Address[243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1147.880 800.000 1148.480 ;
    END
  END Address[243]
  PIN Address[244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1151.960 800.000 1152.560 ;
    END
  END Address[244]
  PIN Address[245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1156.040 800.000 1156.640 ;
    END
  END Address[245]
  PIN Address[246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1160.120 800.000 1160.720 ;
    END
  END Address[246]
  PIN Address[247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1164.200 800.000 1164.800 ;
    END
  END Address[247]
  PIN Address[248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1168.280 800.000 1168.880 ;
    END
  END Address[248]
  PIN Address[249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1172.360 800.000 1172.960 ;
    END
  END Address[249]
  PIN Address[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 254.360 800.000 254.960 ;
    END
  END Address[24]
  PIN Address[250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1176.440 800.000 1177.040 ;
    END
  END Address[250]
  PIN Address[251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1180.520 800.000 1181.120 ;
    END
  END Address[251]
  PIN Address[252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1184.600 800.000 1185.200 ;
    END
  END Address[252]
  PIN Address[253]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1188.680 800.000 1189.280 ;
    END
  END Address[253]
  PIN Address[254]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1192.760 800.000 1193.360 ;
    END
  END Address[254]
  PIN Address[255]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1196.840 800.000 1197.440 ;
    END
  END Address[255]
  PIN Address[256]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1200.920 800.000 1201.520 ;
    END
  END Address[256]
  PIN Address[257]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1205.000 800.000 1205.600 ;
    END
  END Address[257]
  PIN Address[258]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1209.080 800.000 1209.680 ;
    END
  END Address[258]
  PIN Address[259]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1213.160 800.000 1213.760 ;
    END
  END Address[259]
  PIN Address[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 258.440 800.000 259.040 ;
    END
  END Address[25]
  PIN Address[260]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1217.240 800.000 1217.840 ;
    END
  END Address[260]
  PIN Address[261]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1221.320 800.000 1221.920 ;
    END
  END Address[261]
  PIN Address[262]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1225.400 800.000 1226.000 ;
    END
  END Address[262]
  PIN Address[263]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1229.480 800.000 1230.080 ;
    END
  END Address[263]
  PIN Address[264]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1233.560 800.000 1234.160 ;
    END
  END Address[264]
  PIN Address[265]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1237.640 800.000 1238.240 ;
    END
  END Address[265]
  PIN Address[266]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1241.720 800.000 1242.320 ;
    END
  END Address[266]
  PIN Address[267]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1245.800 800.000 1246.400 ;
    END
  END Address[267]
  PIN Address[268]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1249.880 800.000 1250.480 ;
    END
  END Address[268]
  PIN Address[269]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1253.960 800.000 1254.560 ;
    END
  END Address[269]
  PIN Address[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 262.520 800.000 263.120 ;
    END
  END Address[26]
  PIN Address[270]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1258.040 800.000 1258.640 ;
    END
  END Address[270]
  PIN Address[271]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1262.120 800.000 1262.720 ;
    END
  END Address[271]
  PIN Address[272]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1266.200 800.000 1266.800 ;
    END
  END Address[272]
  PIN Address[273]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1270.280 800.000 1270.880 ;
    END
  END Address[273]
  PIN Address[274]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1274.360 800.000 1274.960 ;
    END
  END Address[274]
  PIN Address[275]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1278.440 800.000 1279.040 ;
    END
  END Address[275]
  PIN Address[276]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1282.520 800.000 1283.120 ;
    END
  END Address[276]
  PIN Address[277]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1286.600 800.000 1287.200 ;
    END
  END Address[277]
  PIN Address[278]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1290.680 800.000 1291.280 ;
    END
  END Address[278]
  PIN Address[279]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1294.760 800.000 1295.360 ;
    END
  END Address[279]
  PIN Address[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 266.600 800.000 267.200 ;
    END
  END Address[27]
  PIN Address[280]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1298.840 800.000 1299.440 ;
    END
  END Address[280]
  PIN Address[281]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1302.920 800.000 1303.520 ;
    END
  END Address[281]
  PIN Address[282]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1307.000 800.000 1307.600 ;
    END
  END Address[282]
  PIN Address[283]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1311.080 800.000 1311.680 ;
    END
  END Address[283]
  PIN Address[284]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1315.160 800.000 1315.760 ;
    END
  END Address[284]
  PIN Address[285]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1319.240 800.000 1319.840 ;
    END
  END Address[285]
  PIN Address[286]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1323.320 800.000 1323.920 ;
    END
  END Address[286]
  PIN Address[287]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1327.400 800.000 1328.000 ;
    END
  END Address[287]
  PIN Address[288]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1331.480 800.000 1332.080 ;
    END
  END Address[288]
  PIN Address[289]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1335.560 800.000 1336.160 ;
    END
  END Address[289]
  PIN Address[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 270.680 800.000 271.280 ;
    END
  END Address[28]
  PIN Address[290]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1339.640 800.000 1340.240 ;
    END
  END Address[290]
  PIN Address[291]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1343.720 800.000 1344.320 ;
    END
  END Address[291]
  PIN Address[292]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1347.800 800.000 1348.400 ;
    END
  END Address[292]
  PIN Address[293]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1351.880 800.000 1352.480 ;
    END
  END Address[293]
  PIN Address[294]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1355.960 800.000 1356.560 ;
    END
  END Address[294]
  PIN Address[295]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1360.040 800.000 1360.640 ;
    END
  END Address[295]
  PIN Address[296]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1364.120 800.000 1364.720 ;
    END
  END Address[296]
  PIN Address[297]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1368.200 800.000 1368.800 ;
    END
  END Address[297]
  PIN Address[298]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1372.280 800.000 1372.880 ;
    END
  END Address[298]
  PIN Address[299]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1376.360 800.000 1376.960 ;
    END
  END Address[299]
  PIN Address[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 274.760 800.000 275.360 ;
    END
  END Address[29]
  PIN Address[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 164.600 800.000 165.200 ;
    END
  END Address[2]
  PIN Address[300]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1380.440 800.000 1381.040 ;
    END
  END Address[300]
  PIN Address[301]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1384.520 800.000 1385.120 ;
    END
  END Address[301]
  PIN Address[302]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1388.600 800.000 1389.200 ;
    END
  END Address[302]
  PIN Address[303]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1392.680 800.000 1393.280 ;
    END
  END Address[303]
  PIN Address[304]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1396.760 800.000 1397.360 ;
    END
  END Address[304]
  PIN Address[305]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1400.840 800.000 1401.440 ;
    END
  END Address[305]
  PIN Address[306]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1404.920 800.000 1405.520 ;
    END
  END Address[306]
  PIN Address[307]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1409.000 800.000 1409.600 ;
    END
  END Address[307]
  PIN Address[308]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1413.080 800.000 1413.680 ;
    END
  END Address[308]
  PIN Address[309]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1417.160 800.000 1417.760 ;
    END
  END Address[309]
  PIN Address[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 278.840 800.000 279.440 ;
    END
  END Address[30]
  PIN Address[310]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1421.240 800.000 1421.840 ;
    END
  END Address[310]
  PIN Address[311]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1425.320 800.000 1425.920 ;
    END
  END Address[311]
  PIN Address[312]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1429.400 800.000 1430.000 ;
    END
  END Address[312]
  PIN Address[313]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1433.480 800.000 1434.080 ;
    END
  END Address[313]
  PIN Address[314]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1437.560 800.000 1438.160 ;
    END
  END Address[314]
  PIN Address[315]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1441.640 800.000 1442.240 ;
    END
  END Address[315]
  PIN Address[316]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1445.720 800.000 1446.320 ;
    END
  END Address[316]
  PIN Address[317]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1449.800 800.000 1450.400 ;
    END
  END Address[317]
  PIN Address[318]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1453.880 800.000 1454.480 ;
    END
  END Address[318]
  PIN Address[319]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1457.960 800.000 1458.560 ;
    END
  END Address[319]
  PIN Address[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 282.920 800.000 283.520 ;
    END
  END Address[31]
  PIN Address[320]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1462.040 800.000 1462.640 ;
    END
  END Address[320]
  PIN Address[321]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1466.120 800.000 1466.720 ;
    END
  END Address[321]
  PIN Address[322]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1470.200 800.000 1470.800 ;
    END
  END Address[322]
  PIN Address[323]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1474.280 800.000 1474.880 ;
    END
  END Address[323]
  PIN Address[324]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1478.360 800.000 1478.960 ;
    END
  END Address[324]
  PIN Address[325]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1482.440 800.000 1483.040 ;
    END
  END Address[325]
  PIN Address[326]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1486.520 800.000 1487.120 ;
    END
  END Address[326]
  PIN Address[327]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1490.600 800.000 1491.200 ;
    END
  END Address[327]
  PIN Address[328]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1494.680 800.000 1495.280 ;
    END
  END Address[328]
  PIN Address[329]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1498.760 800.000 1499.360 ;
    END
  END Address[329]
  PIN Address[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 287.000 800.000 287.600 ;
    END
  END Address[32]
  PIN Address[330]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1502.840 800.000 1503.440 ;
    END
  END Address[330]
  PIN Address[331]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1506.920 800.000 1507.520 ;
    END
  END Address[331]
  PIN Address[332]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1511.000 800.000 1511.600 ;
    END
  END Address[332]
  PIN Address[333]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1515.080 800.000 1515.680 ;
    END
  END Address[333]
  PIN Address[334]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1519.160 800.000 1519.760 ;
    END
  END Address[334]
  PIN Address[335]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1523.240 800.000 1523.840 ;
    END
  END Address[335]
  PIN Address[336]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1527.320 800.000 1527.920 ;
    END
  END Address[336]
  PIN Address[337]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1531.400 800.000 1532.000 ;
    END
  END Address[337]
  PIN Address[338]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1535.480 800.000 1536.080 ;
    END
  END Address[338]
  PIN Address[339]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1539.560 800.000 1540.160 ;
    END
  END Address[339]
  PIN Address[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 291.080 800.000 291.680 ;
    END
  END Address[33]
  PIN Address[340]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1543.640 800.000 1544.240 ;
    END
  END Address[340]
  PIN Address[341]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1547.720 800.000 1548.320 ;
    END
  END Address[341]
  PIN Address[342]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1551.800 800.000 1552.400 ;
    END
  END Address[342]
  PIN Address[343]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1555.880 800.000 1556.480 ;
    END
  END Address[343]
  PIN Address[344]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1559.960 800.000 1560.560 ;
    END
  END Address[344]
  PIN Address[345]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1564.040 800.000 1564.640 ;
    END
  END Address[345]
  PIN Address[346]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1568.120 800.000 1568.720 ;
    END
  END Address[346]
  PIN Address[347]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1572.200 800.000 1572.800 ;
    END
  END Address[347]
  PIN Address[348]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1576.280 800.000 1576.880 ;
    END
  END Address[348]
  PIN Address[349]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1580.360 800.000 1580.960 ;
    END
  END Address[349]
  PIN Address[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 295.160 800.000 295.760 ;
    END
  END Address[34]
  PIN Address[350]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1584.440 800.000 1585.040 ;
    END
  END Address[350]
  PIN Address[351]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1588.520 800.000 1589.120 ;
    END
  END Address[351]
  PIN Address[352]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1592.600 800.000 1593.200 ;
    END
  END Address[352]
  PIN Address[353]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1596.680 800.000 1597.280 ;
    END
  END Address[353]
  PIN Address[354]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1600.760 800.000 1601.360 ;
    END
  END Address[354]
  PIN Address[355]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1604.840 800.000 1605.440 ;
    END
  END Address[355]
  PIN Address[356]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1608.920 800.000 1609.520 ;
    END
  END Address[356]
  PIN Address[357]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1613.000 800.000 1613.600 ;
    END
  END Address[357]
  PIN Address[358]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1617.080 800.000 1617.680 ;
    END
  END Address[358]
  PIN Address[359]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1621.160 800.000 1621.760 ;
    END
  END Address[359]
  PIN Address[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 299.240 800.000 299.840 ;
    END
  END Address[35]
  PIN Address[360]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1625.240 800.000 1625.840 ;
    END
  END Address[360]
  PIN Address[361]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1629.320 800.000 1629.920 ;
    END
  END Address[361]
  PIN Address[362]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1633.400 800.000 1634.000 ;
    END
  END Address[362]
  PIN Address[363]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1637.480 800.000 1638.080 ;
    END
  END Address[363]
  PIN Address[364]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1641.560 800.000 1642.160 ;
    END
  END Address[364]
  PIN Address[365]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1645.640 800.000 1646.240 ;
    END
  END Address[365]
  PIN Address[366]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1649.720 800.000 1650.320 ;
    END
  END Address[366]
  PIN Address[367]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1653.800 800.000 1654.400 ;
    END
  END Address[367]
  PIN Address[368]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1657.880 800.000 1658.480 ;
    END
  END Address[368]
  PIN Address[369]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1661.960 800.000 1662.560 ;
    END
  END Address[369]
  PIN Address[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 303.320 800.000 303.920 ;
    END
  END Address[36]
  PIN Address[370]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1666.040 800.000 1666.640 ;
    END
  END Address[370]
  PIN Address[371]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1670.120 800.000 1670.720 ;
    END
  END Address[371]
  PIN Address[372]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1674.200 800.000 1674.800 ;
    END
  END Address[372]
  PIN Address[373]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1678.280 800.000 1678.880 ;
    END
  END Address[373]
  PIN Address[374]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1682.360 800.000 1682.960 ;
    END
  END Address[374]
  PIN Address[375]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1686.440 800.000 1687.040 ;
    END
  END Address[375]
  PIN Address[376]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1690.520 800.000 1691.120 ;
    END
  END Address[376]
  PIN Address[377]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1694.600 800.000 1695.200 ;
    END
  END Address[377]
  PIN Address[378]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1698.680 800.000 1699.280 ;
    END
  END Address[378]
  PIN Address[379]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1702.760 800.000 1703.360 ;
    END
  END Address[379]
  PIN Address[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 307.400 800.000 308.000 ;
    END
  END Address[37]
  PIN Address[380]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1706.840 800.000 1707.440 ;
    END
  END Address[380]
  PIN Address[381]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1710.920 800.000 1711.520 ;
    END
  END Address[381]
  PIN Address[382]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1715.000 800.000 1715.600 ;
    END
  END Address[382]
  PIN Address[383]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1719.080 800.000 1719.680 ;
    END
  END Address[383]
  PIN Address[384]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1723.160 800.000 1723.760 ;
    END
  END Address[384]
  PIN Address[385]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1727.240 800.000 1727.840 ;
    END
  END Address[385]
  PIN Address[386]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1731.320 800.000 1731.920 ;
    END
  END Address[386]
  PIN Address[387]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1735.400 800.000 1736.000 ;
    END
  END Address[387]
  PIN Address[388]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1739.480 800.000 1740.080 ;
    END
  END Address[388]
  PIN Address[389]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1743.560 800.000 1744.160 ;
    END
  END Address[389]
  PIN Address[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 311.480 800.000 312.080 ;
    END
  END Address[38]
  PIN Address[390]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1747.640 800.000 1748.240 ;
    END
  END Address[390]
  PIN Address[391]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1751.720 800.000 1752.320 ;
    END
  END Address[391]
  PIN Address[392]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1755.800 800.000 1756.400 ;
    END
  END Address[392]
  PIN Address[393]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1759.880 800.000 1760.480 ;
    END
  END Address[393]
  PIN Address[394]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1763.960 800.000 1764.560 ;
    END
  END Address[394]
  PIN Address[395]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1768.040 800.000 1768.640 ;
    END
  END Address[395]
  PIN Address[396]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1772.120 800.000 1772.720 ;
    END
  END Address[396]
  PIN Address[397]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1776.200 800.000 1776.800 ;
    END
  END Address[397]
  PIN Address[398]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1780.280 800.000 1780.880 ;
    END
  END Address[398]
  PIN Address[399]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1784.360 800.000 1784.960 ;
    END
  END Address[399]
  PIN Address[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 315.560 800.000 316.160 ;
    END
  END Address[39]
  PIN Address[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 168.680 800.000 169.280 ;
    END
  END Address[3]
  PIN Address[400]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1788.440 800.000 1789.040 ;
    END
  END Address[400]
  PIN Address[401]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1792.520 800.000 1793.120 ;
    END
  END Address[401]
  PIN Address[402]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1796.600 800.000 1797.200 ;
    END
  END Address[402]
  PIN Address[403]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1800.680 800.000 1801.280 ;
    END
  END Address[403]
  PIN Address[404]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1804.760 800.000 1805.360 ;
    END
  END Address[404]
  PIN Address[405]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1808.840 800.000 1809.440 ;
    END
  END Address[405]
  PIN Address[406]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1812.920 800.000 1813.520 ;
    END
  END Address[406]
  PIN Address[407]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1817.000 800.000 1817.600 ;
    END
  END Address[407]
  PIN Address[408]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1821.080 800.000 1821.680 ;
    END
  END Address[408]
  PIN Address[409]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1825.160 800.000 1825.760 ;
    END
  END Address[409]
  PIN Address[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 319.640 800.000 320.240 ;
    END
  END Address[40]
  PIN Address[410]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1829.240 800.000 1829.840 ;
    END
  END Address[410]
  PIN Address[411]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1833.320 800.000 1833.920 ;
    END
  END Address[411]
  PIN Address[412]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1837.400 800.000 1838.000 ;
    END
  END Address[412]
  PIN Address[413]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1841.480 800.000 1842.080 ;
    END
  END Address[413]
  PIN Address[414]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1845.560 800.000 1846.160 ;
    END
  END Address[414]
  PIN Address[415]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1849.640 800.000 1850.240 ;
    END
  END Address[415]
  PIN Address[416]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1853.720 800.000 1854.320 ;
    END
  END Address[416]
  PIN Address[417]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1857.800 800.000 1858.400 ;
    END
  END Address[417]
  PIN Address[418]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1861.880 800.000 1862.480 ;
    END
  END Address[418]
  PIN Address[419]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1865.960 800.000 1866.560 ;
    END
  END Address[419]
  PIN Address[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 323.720 800.000 324.320 ;
    END
  END Address[41]
  PIN Address[420]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1870.040 800.000 1870.640 ;
    END
  END Address[420]
  PIN Address[421]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1874.120 800.000 1874.720 ;
    END
  END Address[421]
  PIN Address[422]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1878.200 800.000 1878.800 ;
    END
  END Address[422]
  PIN Address[423]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1882.280 800.000 1882.880 ;
    END
  END Address[423]
  PIN Address[424]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1886.360 800.000 1886.960 ;
    END
  END Address[424]
  PIN Address[425]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1890.440 800.000 1891.040 ;
    END
  END Address[425]
  PIN Address[426]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1894.520 800.000 1895.120 ;
    END
  END Address[426]
  PIN Address[427]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1898.600 800.000 1899.200 ;
    END
  END Address[427]
  PIN Address[428]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1902.680 800.000 1903.280 ;
    END
  END Address[428]
  PIN Address[429]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1906.760 800.000 1907.360 ;
    END
  END Address[429]
  PIN Address[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 327.800 800.000 328.400 ;
    END
  END Address[42]
  PIN Address[430]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1910.840 800.000 1911.440 ;
    END
  END Address[430]
  PIN Address[431]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1914.920 800.000 1915.520 ;
    END
  END Address[431]
  PIN Address[432]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1919.000 800.000 1919.600 ;
    END
  END Address[432]
  PIN Address[433]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1923.080 800.000 1923.680 ;
    END
  END Address[433]
  PIN Address[434]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1927.160 800.000 1927.760 ;
    END
  END Address[434]
  PIN Address[435]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1931.240 800.000 1931.840 ;
    END
  END Address[435]
  PIN Address[436]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1935.320 800.000 1935.920 ;
    END
  END Address[436]
  PIN Address[437]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1939.400 800.000 1940.000 ;
    END
  END Address[437]
  PIN Address[438]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1943.480 800.000 1944.080 ;
    END
  END Address[438]
  PIN Address[439]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1947.560 800.000 1948.160 ;
    END
  END Address[439]
  PIN Address[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 331.880 800.000 332.480 ;
    END
  END Address[43]
  PIN Address[440]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1951.640 800.000 1952.240 ;
    END
  END Address[440]
  PIN Address[441]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1955.720 800.000 1956.320 ;
    END
  END Address[441]
  PIN Address[442]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1959.800 800.000 1960.400 ;
    END
  END Address[442]
  PIN Address[443]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1963.880 800.000 1964.480 ;
    END
  END Address[443]
  PIN Address[444]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1967.960 800.000 1968.560 ;
    END
  END Address[444]
  PIN Address[445]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1972.040 800.000 1972.640 ;
    END
  END Address[445]
  PIN Address[446]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1976.120 800.000 1976.720 ;
    END
  END Address[446]
  PIN Address[447]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1980.200 800.000 1980.800 ;
    END
  END Address[447]
  PIN Address[448]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1984.280 800.000 1984.880 ;
    END
  END Address[448]
  PIN Address[449]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1988.360 800.000 1988.960 ;
    END
  END Address[449]
  PIN Address[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 335.960 800.000 336.560 ;
    END
  END Address[44]
  PIN Address[450]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1992.440 800.000 1993.040 ;
    END
  END Address[450]
  PIN Address[451]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 1996.520 800.000 1997.120 ;
    END
  END Address[451]
  PIN Address[452]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 2000.600 800.000 2001.200 ;
    END
  END Address[452]
  PIN Address[453]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 2004.680 800.000 2005.280 ;
    END
  END Address[453]
  PIN Address[454]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 2008.760 800.000 2009.360 ;
    END
  END Address[454]
  PIN Address[455]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 2012.840 800.000 2013.440 ;
    END
  END Address[455]
  PIN Address[456]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 2016.920 800.000 2017.520 ;
    END
  END Address[456]
  PIN Address[457]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 2021.000 800.000 2021.600 ;
    END
  END Address[457]
  PIN Address[458]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 2025.080 800.000 2025.680 ;
    END
  END Address[458]
  PIN Address[459]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 2029.160 800.000 2029.760 ;
    END
  END Address[459]
  PIN Address[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 340.040 800.000 340.640 ;
    END
  END Address[45]
  PIN Address[460]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 2033.240 800.000 2033.840 ;
    END
  END Address[460]
  PIN Address[461]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 2037.320 800.000 2037.920 ;
    END
  END Address[461]
  PIN Address[462]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 2041.400 800.000 2042.000 ;
    END
  END Address[462]
  PIN Address[463]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 2045.480 800.000 2046.080 ;
    END
  END Address[463]
  PIN Address[464]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 2049.560 800.000 2050.160 ;
    END
  END Address[464]
  PIN Address[465]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 2053.640 800.000 2054.240 ;
    END
  END Address[465]
  PIN Address[466]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 2057.720 800.000 2058.320 ;
    END
  END Address[466]
  PIN Address[467]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 2061.800 800.000 2062.400 ;
    END
  END Address[467]
  PIN Address[468]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 2065.880 800.000 2066.480 ;
    END
  END Address[468]
  PIN Address[469]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 2069.960 800.000 2070.560 ;
    END
  END Address[469]
  PIN Address[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 344.120 800.000 344.720 ;
    END
  END Address[46]
  PIN Address[470]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 2074.040 800.000 2074.640 ;
    END
  END Address[470]
  PIN Address[471]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 2078.120 800.000 2078.720 ;
    END
  END Address[471]
  PIN Address[472]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 2082.200 800.000 2082.800 ;
    END
  END Address[472]
  PIN Address[473]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 2086.280 800.000 2086.880 ;
    END
  END Address[473]
  PIN Address[474]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 2090.360 800.000 2090.960 ;
    END
  END Address[474]
  PIN Address[475]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 2094.440 800.000 2095.040 ;
    END
  END Address[475]
  PIN Address[476]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 2098.520 800.000 2099.120 ;
    END
  END Address[476]
  PIN Address[477]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 2102.600 800.000 2103.200 ;
    END
  END Address[477]
  PIN Address[478]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 2106.680 800.000 2107.280 ;
    END
  END Address[478]
  PIN Address[479]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 796.000 2110.760 800.000 2111.360 ;
    END
  END Address[479]
  PIN Address[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 348.200 800.000 348.800 ;
    END
  END Address[47]
  PIN Address[480]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 2114.840 800.000 2115.440 ;
    END
  END Address[480]
  PIN Address[481]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 2118.920 800.000 2119.520 ;
    END
  END Address[481]
  PIN Address[482]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 2123.000 800.000 2123.600 ;
    END
  END Address[482]
  PIN Address[483]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 2127.080 800.000 2127.680 ;
    END
  END Address[483]
  PIN Address[484]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 2131.160 800.000 2131.760 ;
    END
  END Address[484]
  PIN Address[485]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 2135.240 800.000 2135.840 ;
    END
  END Address[485]
  PIN Address[486]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 2139.320 800.000 2139.920 ;
    END
  END Address[486]
  PIN Address[487]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 2143.400 800.000 2144.000 ;
    END
  END Address[487]
  PIN Address[488]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 2147.480 800.000 2148.080 ;
    END
  END Address[488]
  PIN Address[489]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 2151.560 800.000 2152.160 ;
    END
  END Address[489]
  PIN Address[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 352.280 800.000 352.880 ;
    END
  END Address[48]
  PIN Address[490]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 2155.640 800.000 2156.240 ;
    END
  END Address[490]
  PIN Address[491]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 2159.720 800.000 2160.320 ;
    END
  END Address[491]
  PIN Address[492]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 2163.800 800.000 2164.400 ;
    END
  END Address[492]
  PIN Address[493]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 2167.880 800.000 2168.480 ;
    END
  END Address[493]
  PIN Address[494]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 2171.960 800.000 2172.560 ;
    END
  END Address[494]
  PIN Address[495]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 2176.040 800.000 2176.640 ;
    END
  END Address[495]
  PIN Address[496]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 2180.120 800.000 2180.720 ;
    END
  END Address[496]
  PIN Address[497]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 2184.200 800.000 2184.800 ;
    END
  END Address[497]
  PIN Address[498]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 2188.280 800.000 2188.880 ;
    END
  END Address[498]
  PIN Address[499]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 2192.360 800.000 2192.960 ;
    END
  END Address[499]
  PIN Address[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 356.360 800.000 356.960 ;
    END
  END Address[49]
  PIN Address[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 172.760 800.000 173.360 ;
    END
  END Address[4]
  PIN Address[500]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 2196.440 800.000 2197.040 ;
    END
  END Address[500]
  PIN Address[501]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 2200.520 800.000 2201.120 ;
    END
  END Address[501]
  PIN Address[502]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 2204.600 800.000 2205.200 ;
    END
  END Address[502]
  PIN Address[503]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 2208.680 800.000 2209.280 ;
    END
  END Address[503]
  PIN Address[504]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 2212.760 800.000 2213.360 ;
    END
  END Address[504]
  PIN Address[505]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 2216.840 800.000 2217.440 ;
    END
  END Address[505]
  PIN Address[506]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 2220.920 800.000 2221.520 ;
    END
  END Address[506]
  PIN Address[507]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 2225.000 800.000 2225.600 ;
    END
  END Address[507]
  PIN Address[508]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 2229.080 800.000 2229.680 ;
    END
  END Address[508]
  PIN Address[509]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 2233.160 800.000 2233.760 ;
    END
  END Address[509]
  PIN Address[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 360.440 800.000 361.040 ;
    END
  END Address[50]
  PIN Address[510]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 2237.240 800.000 2237.840 ;
    END
  END Address[510]
  PIN Address[511]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 2241.320 800.000 2241.920 ;
    END
  END Address[511]
  PIN Address[512]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 156.440 4.000 157.040 ;
    END
  END Address[512]
  PIN Address[513]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 160.520 4.000 161.120 ;
    END
  END Address[513]
  PIN Address[514]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 164.600 4.000 165.200 ;
    END
  END Address[514]
  PIN Address[515]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.680 4.000 169.280 ;
    END
  END Address[515]
  PIN Address[516]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.760 4.000 173.360 ;
    END
  END Address[516]
  PIN Address[517]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END Address[517]
  PIN Address[518]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.920 4.000 181.520 ;
    END
  END Address[518]
  PIN Address[519]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.000 4.000 185.600 ;
    END
  END Address[519]
  PIN Address[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 364.520 800.000 365.120 ;
    END
  END Address[51]
  PIN Address[520]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.080 4.000 189.680 ;
    END
  END Address[520]
  PIN Address[521]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.160 4.000 193.760 ;
    END
  END Address[521]
  PIN Address[522]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.240 4.000 197.840 ;
    END
  END Address[522]
  PIN Address[523]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 201.320 4.000 201.920 ;
    END
  END Address[523]
  PIN Address[524]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 205.400 4.000 206.000 ;
    END
  END Address[524]
  PIN Address[525]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 209.480 4.000 210.080 ;
    END
  END Address[525]
  PIN Address[526]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 213.560 4.000 214.160 ;
    END
  END Address[526]
  PIN Address[527]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END Address[527]
  PIN Address[528]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.720 4.000 222.320 ;
    END
  END Address[528]
  PIN Address[529]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.800 4.000 226.400 ;
    END
  END Address[529]
  PIN Address[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 368.600 800.000 369.200 ;
    END
  END Address[52]
  PIN Address[530]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.880 4.000 230.480 ;
    END
  END Address[530]
  PIN Address[531]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 233.960 4.000 234.560 ;
    END
  END Address[531]
  PIN Address[532]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.040 4.000 238.640 ;
    END
  END Address[532]
  PIN Address[533]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 242.120 4.000 242.720 ;
    END
  END Address[533]
  PIN Address[534]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 246.200 4.000 246.800 ;
    END
  END Address[534]
  PIN Address[535]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 250.280 4.000 250.880 ;
    END
  END Address[535]
  PIN Address[536]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 254.360 4.000 254.960 ;
    END
  END Address[536]
  PIN Address[537]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END Address[537]
  PIN Address[538]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 262.520 4.000 263.120 ;
    END
  END Address[538]
  PIN Address[539]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 266.600 4.000 267.200 ;
    END
  END Address[539]
  PIN Address[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 372.680 800.000 373.280 ;
    END
  END Address[53]
  PIN Address[540]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.680 4.000 271.280 ;
    END
  END Address[540]
  PIN Address[541]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 274.760 4.000 275.360 ;
    END
  END Address[541]
  PIN Address[542]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.840 4.000 279.440 ;
    END
  END Address[542]
  PIN Address[543]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.920 4.000 283.520 ;
    END
  END Address[543]
  PIN Address[544]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 287.000 4.000 287.600 ;
    END
  END Address[544]
  PIN Address[545]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 291.080 4.000 291.680 ;
    END
  END Address[545]
  PIN Address[546]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.160 4.000 295.760 ;
    END
  END Address[546]
  PIN Address[547]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END Address[547]
  PIN Address[548]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 303.320 4.000 303.920 ;
    END
  END Address[548]
  PIN Address[549]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 307.400 4.000 308.000 ;
    END
  END Address[549]
  PIN Address[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 376.760 800.000 377.360 ;
    END
  END Address[54]
  PIN Address[550]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 311.480 4.000 312.080 ;
    END
  END Address[550]
  PIN Address[551]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 315.560 4.000 316.160 ;
    END
  END Address[551]
  PIN Address[552]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 319.640 4.000 320.240 ;
    END
  END Address[552]
  PIN Address[553]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.720 4.000 324.320 ;
    END
  END Address[553]
  PIN Address[554]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 327.800 4.000 328.400 ;
    END
  END Address[554]
  PIN Address[555]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 331.880 4.000 332.480 ;
    END
  END Address[555]
  PIN Address[556]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 335.960 4.000 336.560 ;
    END
  END Address[556]
  PIN Address[557]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.040 4.000 340.640 ;
    END
  END Address[557]
  PIN Address[558]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 344.120 4.000 344.720 ;
    END
  END Address[558]
  PIN Address[559]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 348.200 4.000 348.800 ;
    END
  END Address[559]
  PIN Address[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 380.840 800.000 381.440 ;
    END
  END Address[55]
  PIN Address[560]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 352.280 4.000 352.880 ;
    END
  END Address[560]
  PIN Address[561]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 356.360 4.000 356.960 ;
    END
  END Address[561]
  PIN Address[562]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 360.440 4.000 361.040 ;
    END
  END Address[562]
  PIN Address[563]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 364.520 4.000 365.120 ;
    END
  END Address[563]
  PIN Address[564]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 368.600 4.000 369.200 ;
    END
  END Address[564]
  PIN Address[565]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 372.680 4.000 373.280 ;
    END
  END Address[565]
  PIN Address[566]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 376.760 4.000 377.360 ;
    END
  END Address[566]
  PIN Address[567]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 4.000 381.440 ;
    END
  END Address[567]
  PIN Address[568]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.920 4.000 385.520 ;
    END
  END Address[568]
  PIN Address[569]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 389.000 4.000 389.600 ;
    END
  END Address[569]
  PIN Address[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 384.920 800.000 385.520 ;
    END
  END Address[56]
  PIN Address[570]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 393.080 4.000 393.680 ;
    END
  END Address[570]
  PIN Address[571]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.160 4.000 397.760 ;
    END
  END Address[571]
  PIN Address[572]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 401.240 4.000 401.840 ;
    END
  END Address[572]
  PIN Address[573]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 405.320 4.000 405.920 ;
    END
  END Address[573]
  PIN Address[574]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 409.400 4.000 410.000 ;
    END
  END Address[574]
  PIN Address[575]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 413.480 4.000 414.080 ;
    END
  END Address[575]
  PIN Address[576]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 417.560 4.000 418.160 ;
    END
  END Address[576]
  PIN Address[577]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 421.640 4.000 422.240 ;
    END
  END Address[577]
  PIN Address[578]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 425.720 4.000 426.320 ;
    END
  END Address[578]
  PIN Address[579]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 429.800 4.000 430.400 ;
    END
  END Address[579]
  PIN Address[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 389.000 800.000 389.600 ;
    END
  END Address[57]
  PIN Address[580]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 433.880 4.000 434.480 ;
    END
  END Address[580]
  PIN Address[581]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 437.960 4.000 438.560 ;
    END
  END Address[581]
  PIN Address[582]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 442.040 4.000 442.640 ;
    END
  END Address[582]
  PIN Address[583]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 446.120 4.000 446.720 ;
    END
  END Address[583]
  PIN Address[584]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 450.200 4.000 450.800 ;
    END
  END Address[584]
  PIN Address[585]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 454.280 4.000 454.880 ;
    END
  END Address[585]
  PIN Address[586]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 458.360 4.000 458.960 ;
    END
  END Address[586]
  PIN Address[587]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 462.440 4.000 463.040 ;
    END
  END Address[587]
  PIN Address[588]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 466.520 4.000 467.120 ;
    END
  END Address[588]
  PIN Address[589]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 470.600 4.000 471.200 ;
    END
  END Address[589]
  PIN Address[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 393.080 800.000 393.680 ;
    END
  END Address[58]
  PIN Address[590]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 474.680 4.000 475.280 ;
    END
  END Address[590]
  PIN Address[591]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 478.760 4.000 479.360 ;
    END
  END Address[591]
  PIN Address[592]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 482.840 4.000 483.440 ;
    END
  END Address[592]
  PIN Address[593]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 486.920 4.000 487.520 ;
    END
  END Address[593]
  PIN Address[594]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 491.000 4.000 491.600 ;
    END
  END Address[594]
  PIN Address[595]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 495.080 4.000 495.680 ;
    END
  END Address[595]
  PIN Address[596]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 499.160 4.000 499.760 ;
    END
  END Address[596]
  PIN Address[597]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 503.240 4.000 503.840 ;
    END
  END Address[597]
  PIN Address[598]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 507.320 4.000 507.920 ;
    END
  END Address[598]
  PIN Address[599]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 511.400 4.000 512.000 ;
    END
  END Address[599]
  PIN Address[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 397.160 800.000 397.760 ;
    END
  END Address[59]
  PIN Address[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 176.840 800.000 177.440 ;
    END
  END Address[5]
  PIN Address[600]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 515.480 4.000 516.080 ;
    END
  END Address[600]
  PIN Address[601]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 519.560 4.000 520.160 ;
    END
  END Address[601]
  PIN Address[602]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 523.640 4.000 524.240 ;
    END
  END Address[602]
  PIN Address[603]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 527.720 4.000 528.320 ;
    END
  END Address[603]
  PIN Address[604]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 531.800 4.000 532.400 ;
    END
  END Address[604]
  PIN Address[605]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 535.880 4.000 536.480 ;
    END
  END Address[605]
  PIN Address[606]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 539.960 4.000 540.560 ;
    END
  END Address[606]
  PIN Address[607]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 544.040 4.000 544.640 ;
    END
  END Address[607]
  PIN Address[608]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 548.120 4.000 548.720 ;
    END
  END Address[608]
  PIN Address[609]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 552.200 4.000 552.800 ;
    END
  END Address[609]
  PIN Address[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 401.240 800.000 401.840 ;
    END
  END Address[60]
  PIN Address[610]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 556.280 4.000 556.880 ;
    END
  END Address[610]
  PIN Address[611]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 560.360 4.000 560.960 ;
    END
  END Address[611]
  PIN Address[612]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 564.440 4.000 565.040 ;
    END
  END Address[612]
  PIN Address[613]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 568.520 4.000 569.120 ;
    END
  END Address[613]
  PIN Address[614]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 572.600 4.000 573.200 ;
    END
  END Address[614]
  PIN Address[615]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 576.680 4.000 577.280 ;
    END
  END Address[615]
  PIN Address[616]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 580.760 4.000 581.360 ;
    END
  END Address[616]
  PIN Address[617]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 584.840 4.000 585.440 ;
    END
  END Address[617]
  PIN Address[618]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 588.920 4.000 589.520 ;
    END
  END Address[618]
  PIN Address[619]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 593.000 4.000 593.600 ;
    END
  END Address[619]
  PIN Address[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 405.320 800.000 405.920 ;
    END
  END Address[61]
  PIN Address[620]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 597.080 4.000 597.680 ;
    END
  END Address[620]
  PIN Address[621]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 601.160 4.000 601.760 ;
    END
  END Address[621]
  PIN Address[622]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 605.240 4.000 605.840 ;
    END
  END Address[622]
  PIN Address[623]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 609.320 4.000 609.920 ;
    END
  END Address[623]
  PIN Address[624]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 613.400 4.000 614.000 ;
    END
  END Address[624]
  PIN Address[625]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 617.480 4.000 618.080 ;
    END
  END Address[625]
  PIN Address[626]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 621.560 4.000 622.160 ;
    END
  END Address[626]
  PIN Address[627]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 625.640 4.000 626.240 ;
    END
  END Address[627]
  PIN Address[628]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 629.720 4.000 630.320 ;
    END
  END Address[628]
  PIN Address[629]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 633.800 4.000 634.400 ;
    END
  END Address[629]
  PIN Address[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 409.400 800.000 410.000 ;
    END
  END Address[62]
  PIN Address[630]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 637.880 4.000 638.480 ;
    END
  END Address[630]
  PIN Address[631]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 641.960 4.000 642.560 ;
    END
  END Address[631]
  PIN Address[632]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 646.040 4.000 646.640 ;
    END
  END Address[632]
  PIN Address[633]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 650.120 4.000 650.720 ;
    END
  END Address[633]
  PIN Address[634]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 654.200 4.000 654.800 ;
    END
  END Address[634]
  PIN Address[635]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 658.280 4.000 658.880 ;
    END
  END Address[635]
  PIN Address[636]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 662.360 4.000 662.960 ;
    END
  END Address[636]
  PIN Address[637]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 666.440 4.000 667.040 ;
    END
  END Address[637]
  PIN Address[638]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 670.520 4.000 671.120 ;
    END
  END Address[638]
  PIN Address[639]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 674.600 4.000 675.200 ;
    END
  END Address[639]
  PIN Address[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 413.480 800.000 414.080 ;
    END
  END Address[63]
  PIN Address[640]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 678.680 4.000 679.280 ;
    END
  END Address[640]
  PIN Address[641]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 682.760 4.000 683.360 ;
    END
  END Address[641]
  PIN Address[642]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 686.840 4.000 687.440 ;
    END
  END Address[642]
  PIN Address[643]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 690.920 4.000 691.520 ;
    END
  END Address[643]
  PIN Address[644]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 695.000 4.000 695.600 ;
    END
  END Address[644]
  PIN Address[645]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 699.080 4.000 699.680 ;
    END
  END Address[645]
  PIN Address[646]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 703.160 4.000 703.760 ;
    END
  END Address[646]
  PIN Address[647]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 707.240 4.000 707.840 ;
    END
  END Address[647]
  PIN Address[648]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 711.320 4.000 711.920 ;
    END
  END Address[648]
  PIN Address[649]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 715.400 4.000 716.000 ;
    END
  END Address[649]
  PIN Address[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 417.560 800.000 418.160 ;
    END
  END Address[64]
  PIN Address[650]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 719.480 4.000 720.080 ;
    END
  END Address[650]
  PIN Address[651]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 723.560 4.000 724.160 ;
    END
  END Address[651]
  PIN Address[652]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 727.640 4.000 728.240 ;
    END
  END Address[652]
  PIN Address[653]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 731.720 4.000 732.320 ;
    END
  END Address[653]
  PIN Address[654]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 735.800 4.000 736.400 ;
    END
  END Address[654]
  PIN Address[655]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 739.880 4.000 740.480 ;
    END
  END Address[655]
  PIN Address[656]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 743.960 4.000 744.560 ;
    END
  END Address[656]
  PIN Address[657]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 748.040 4.000 748.640 ;
    END
  END Address[657]
  PIN Address[658]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 752.120 4.000 752.720 ;
    END
  END Address[658]
  PIN Address[659]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 756.200 4.000 756.800 ;
    END
  END Address[659]
  PIN Address[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 421.640 800.000 422.240 ;
    END
  END Address[65]
  PIN Address[660]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 760.280 4.000 760.880 ;
    END
  END Address[660]
  PIN Address[661]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 764.360 4.000 764.960 ;
    END
  END Address[661]
  PIN Address[662]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 768.440 4.000 769.040 ;
    END
  END Address[662]
  PIN Address[663]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 772.520 4.000 773.120 ;
    END
  END Address[663]
  PIN Address[664]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 776.600 4.000 777.200 ;
    END
  END Address[664]
  PIN Address[665]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 780.680 4.000 781.280 ;
    END
  END Address[665]
  PIN Address[666]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 784.760 4.000 785.360 ;
    END
  END Address[666]
  PIN Address[667]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 788.840 4.000 789.440 ;
    END
  END Address[667]
  PIN Address[668]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 792.920 4.000 793.520 ;
    END
  END Address[668]
  PIN Address[669]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 797.000 4.000 797.600 ;
    END
  END Address[669]
  PIN Address[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 425.720 800.000 426.320 ;
    END
  END Address[66]
  PIN Address[670]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 801.080 4.000 801.680 ;
    END
  END Address[670]
  PIN Address[671]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 805.160 4.000 805.760 ;
    END
  END Address[671]
  PIN Address[672]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 809.240 4.000 809.840 ;
    END
  END Address[672]
  PIN Address[673]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 813.320 4.000 813.920 ;
    END
  END Address[673]
  PIN Address[674]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 817.400 4.000 818.000 ;
    END
  END Address[674]
  PIN Address[675]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 821.480 4.000 822.080 ;
    END
  END Address[675]
  PIN Address[676]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 825.560 4.000 826.160 ;
    END
  END Address[676]
  PIN Address[677]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 829.640 4.000 830.240 ;
    END
  END Address[677]
  PIN Address[678]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 833.720 4.000 834.320 ;
    END
  END Address[678]
  PIN Address[679]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 837.800 4.000 838.400 ;
    END
  END Address[679]
  PIN Address[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 429.800 800.000 430.400 ;
    END
  END Address[67]
  PIN Address[680]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 841.880 4.000 842.480 ;
    END
  END Address[680]
  PIN Address[681]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 845.960 4.000 846.560 ;
    END
  END Address[681]
  PIN Address[682]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 850.040 4.000 850.640 ;
    END
  END Address[682]
  PIN Address[683]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 854.120 4.000 854.720 ;
    END
  END Address[683]
  PIN Address[684]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 858.200 4.000 858.800 ;
    END
  END Address[684]
  PIN Address[685]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 862.280 4.000 862.880 ;
    END
  END Address[685]
  PIN Address[686]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 866.360 4.000 866.960 ;
    END
  END Address[686]
  PIN Address[687]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 870.440 4.000 871.040 ;
    END
  END Address[687]
  PIN Address[688]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 874.520 4.000 875.120 ;
    END
  END Address[688]
  PIN Address[689]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 878.600 4.000 879.200 ;
    END
  END Address[689]
  PIN Address[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 433.880 800.000 434.480 ;
    END
  END Address[68]
  PIN Address[690]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 882.680 4.000 883.280 ;
    END
  END Address[690]
  PIN Address[691]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 886.760 4.000 887.360 ;
    END
  END Address[691]
  PIN Address[692]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 890.840 4.000 891.440 ;
    END
  END Address[692]
  PIN Address[693]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 894.920 4.000 895.520 ;
    END
  END Address[693]
  PIN Address[694]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 899.000 4.000 899.600 ;
    END
  END Address[694]
  PIN Address[695]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 903.080 4.000 903.680 ;
    END
  END Address[695]
  PIN Address[696]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 907.160 4.000 907.760 ;
    END
  END Address[696]
  PIN Address[697]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 911.240 4.000 911.840 ;
    END
  END Address[697]
  PIN Address[698]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 915.320 4.000 915.920 ;
    END
  END Address[698]
  PIN Address[699]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 919.400 4.000 920.000 ;
    END
  END Address[699]
  PIN Address[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 437.960 800.000 438.560 ;
    END
  END Address[69]
  PIN Address[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 180.920 800.000 181.520 ;
    END
  END Address[6]
  PIN Address[700]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 923.480 4.000 924.080 ;
    END
  END Address[700]
  PIN Address[701]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 927.560 4.000 928.160 ;
    END
  END Address[701]
  PIN Address[702]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 931.640 4.000 932.240 ;
    END
  END Address[702]
  PIN Address[703]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 935.720 4.000 936.320 ;
    END
  END Address[703]
  PIN Address[704]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 939.800 4.000 940.400 ;
    END
  END Address[704]
  PIN Address[705]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 943.880 4.000 944.480 ;
    END
  END Address[705]
  PIN Address[706]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 947.960 4.000 948.560 ;
    END
  END Address[706]
  PIN Address[707]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 952.040 4.000 952.640 ;
    END
  END Address[707]
  PIN Address[708]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 956.120 4.000 956.720 ;
    END
  END Address[708]
  PIN Address[709]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 960.200 4.000 960.800 ;
    END
  END Address[709]
  PIN Address[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 442.040 800.000 442.640 ;
    END
  END Address[70]
  PIN Address[710]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 964.280 4.000 964.880 ;
    END
  END Address[710]
  PIN Address[711]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 968.360 4.000 968.960 ;
    END
  END Address[711]
  PIN Address[712]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 972.440 4.000 973.040 ;
    END
  END Address[712]
  PIN Address[713]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 976.520 4.000 977.120 ;
    END
  END Address[713]
  PIN Address[714]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 980.600 4.000 981.200 ;
    END
  END Address[714]
  PIN Address[715]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 984.680 4.000 985.280 ;
    END
  END Address[715]
  PIN Address[716]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 988.760 4.000 989.360 ;
    END
  END Address[716]
  PIN Address[717]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 992.840 4.000 993.440 ;
    END
  END Address[717]
  PIN Address[718]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 996.920 4.000 997.520 ;
    END
  END Address[718]
  PIN Address[719]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1001.000 4.000 1001.600 ;
    END
  END Address[719]
  PIN Address[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 446.120 800.000 446.720 ;
    END
  END Address[71]
  PIN Address[720]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1005.080 4.000 1005.680 ;
    END
  END Address[720]
  PIN Address[721]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1009.160 4.000 1009.760 ;
    END
  END Address[721]
  PIN Address[722]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1013.240 4.000 1013.840 ;
    END
  END Address[722]
  PIN Address[723]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1017.320 4.000 1017.920 ;
    END
  END Address[723]
  PIN Address[724]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1021.400 4.000 1022.000 ;
    END
  END Address[724]
  PIN Address[725]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1025.480 4.000 1026.080 ;
    END
  END Address[725]
  PIN Address[726]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1029.560 4.000 1030.160 ;
    END
  END Address[726]
  PIN Address[727]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1033.640 4.000 1034.240 ;
    END
  END Address[727]
  PIN Address[728]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1037.720 4.000 1038.320 ;
    END
  END Address[728]
  PIN Address[729]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1041.800 4.000 1042.400 ;
    END
  END Address[729]
  PIN Address[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 450.200 800.000 450.800 ;
    END
  END Address[72]
  PIN Address[730]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1045.880 4.000 1046.480 ;
    END
  END Address[730]
  PIN Address[731]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1049.960 4.000 1050.560 ;
    END
  END Address[731]
  PIN Address[732]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1054.040 4.000 1054.640 ;
    END
  END Address[732]
  PIN Address[733]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1058.120 4.000 1058.720 ;
    END
  END Address[733]
  PIN Address[734]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1062.200 4.000 1062.800 ;
    END
  END Address[734]
  PIN Address[735]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1066.280 4.000 1066.880 ;
    END
  END Address[735]
  PIN Address[736]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1070.360 4.000 1070.960 ;
    END
  END Address[736]
  PIN Address[737]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1074.440 4.000 1075.040 ;
    END
  END Address[737]
  PIN Address[738]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1078.520 4.000 1079.120 ;
    END
  END Address[738]
  PIN Address[739]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1082.600 4.000 1083.200 ;
    END
  END Address[739]
  PIN Address[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 454.280 800.000 454.880 ;
    END
  END Address[73]
  PIN Address[740]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1086.680 4.000 1087.280 ;
    END
  END Address[740]
  PIN Address[741]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1090.760 4.000 1091.360 ;
    END
  END Address[741]
  PIN Address[742]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1094.840 4.000 1095.440 ;
    END
  END Address[742]
  PIN Address[743]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1098.920 4.000 1099.520 ;
    END
  END Address[743]
  PIN Address[744]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1103.000 4.000 1103.600 ;
    END
  END Address[744]
  PIN Address[745]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1107.080 4.000 1107.680 ;
    END
  END Address[745]
  PIN Address[746]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1111.160 4.000 1111.760 ;
    END
  END Address[746]
  PIN Address[747]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1115.240 4.000 1115.840 ;
    END
  END Address[747]
  PIN Address[748]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1119.320 4.000 1119.920 ;
    END
  END Address[748]
  PIN Address[749]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1123.400 4.000 1124.000 ;
    END
  END Address[749]
  PIN Address[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 458.360 800.000 458.960 ;
    END
  END Address[74]
  PIN Address[750]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1127.480 4.000 1128.080 ;
    END
  END Address[750]
  PIN Address[751]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1131.560 4.000 1132.160 ;
    END
  END Address[751]
  PIN Address[752]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1135.640 4.000 1136.240 ;
    END
  END Address[752]
  PIN Address[753]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1139.720 4.000 1140.320 ;
    END
  END Address[753]
  PIN Address[754]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1143.800 4.000 1144.400 ;
    END
  END Address[754]
  PIN Address[755]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1147.880 4.000 1148.480 ;
    END
  END Address[755]
  PIN Address[756]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1151.960 4.000 1152.560 ;
    END
  END Address[756]
  PIN Address[757]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1156.040 4.000 1156.640 ;
    END
  END Address[757]
  PIN Address[758]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1160.120 4.000 1160.720 ;
    END
  END Address[758]
  PIN Address[759]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1164.200 4.000 1164.800 ;
    END
  END Address[759]
  PIN Address[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 462.440 800.000 463.040 ;
    END
  END Address[75]
  PIN Address[760]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1168.280 4.000 1168.880 ;
    END
  END Address[760]
  PIN Address[761]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1172.360 4.000 1172.960 ;
    END
  END Address[761]
  PIN Address[762]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1176.440 4.000 1177.040 ;
    END
  END Address[762]
  PIN Address[763]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1180.520 4.000 1181.120 ;
    END
  END Address[763]
  PIN Address[764]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1184.600 4.000 1185.200 ;
    END
  END Address[764]
  PIN Address[765]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1188.680 4.000 1189.280 ;
    END
  END Address[765]
  PIN Address[766]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1192.760 4.000 1193.360 ;
    END
  END Address[766]
  PIN Address[767]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1196.840 4.000 1197.440 ;
    END
  END Address[767]
  PIN Address[768]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1200.920 4.000 1201.520 ;
    END
  END Address[768]
  PIN Address[769]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1205.000 4.000 1205.600 ;
    END
  END Address[769]
  PIN Address[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 466.520 800.000 467.120 ;
    END
  END Address[76]
  PIN Address[770]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1209.080 4.000 1209.680 ;
    END
  END Address[770]
  PIN Address[771]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1213.160 4.000 1213.760 ;
    END
  END Address[771]
  PIN Address[772]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1217.240 4.000 1217.840 ;
    END
  END Address[772]
  PIN Address[773]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1221.320 4.000 1221.920 ;
    END
  END Address[773]
  PIN Address[774]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1225.400 4.000 1226.000 ;
    END
  END Address[774]
  PIN Address[775]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1229.480 4.000 1230.080 ;
    END
  END Address[775]
  PIN Address[776]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1233.560 4.000 1234.160 ;
    END
  END Address[776]
  PIN Address[777]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1237.640 4.000 1238.240 ;
    END
  END Address[777]
  PIN Address[778]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1241.720 4.000 1242.320 ;
    END
  END Address[778]
  PIN Address[779]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1245.800 4.000 1246.400 ;
    END
  END Address[779]
  PIN Address[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 470.600 800.000 471.200 ;
    END
  END Address[77]
  PIN Address[780]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1249.880 4.000 1250.480 ;
    END
  END Address[780]
  PIN Address[781]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1253.960 4.000 1254.560 ;
    END
  END Address[781]
  PIN Address[782]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1258.040 4.000 1258.640 ;
    END
  END Address[782]
  PIN Address[783]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1262.120 4.000 1262.720 ;
    END
  END Address[783]
  PIN Address[784]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1266.200 4.000 1266.800 ;
    END
  END Address[784]
  PIN Address[785]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1270.280 4.000 1270.880 ;
    END
  END Address[785]
  PIN Address[786]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1274.360 4.000 1274.960 ;
    END
  END Address[786]
  PIN Address[787]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1278.440 4.000 1279.040 ;
    END
  END Address[787]
  PIN Address[788]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1282.520 4.000 1283.120 ;
    END
  END Address[788]
  PIN Address[789]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1286.600 4.000 1287.200 ;
    END
  END Address[789]
  PIN Address[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 474.680 800.000 475.280 ;
    END
  END Address[78]
  PIN Address[790]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1290.680 4.000 1291.280 ;
    END
  END Address[790]
  PIN Address[791]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1294.760 4.000 1295.360 ;
    END
  END Address[791]
  PIN Address[792]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1298.840 4.000 1299.440 ;
    END
  END Address[792]
  PIN Address[793]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1302.920 4.000 1303.520 ;
    END
  END Address[793]
  PIN Address[794]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1307.000 4.000 1307.600 ;
    END
  END Address[794]
  PIN Address[795]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1311.080 4.000 1311.680 ;
    END
  END Address[795]
  PIN Address[796]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1315.160 4.000 1315.760 ;
    END
  END Address[796]
  PIN Address[797]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1319.240 4.000 1319.840 ;
    END
  END Address[797]
  PIN Address[798]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1323.320 4.000 1323.920 ;
    END
  END Address[798]
  PIN Address[799]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1327.400 4.000 1328.000 ;
    END
  END Address[799]
  PIN Address[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 478.760 800.000 479.360 ;
    END
  END Address[79]
  PIN Address[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 185.000 800.000 185.600 ;
    END
  END Address[7]
  PIN Address[800]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1331.480 4.000 1332.080 ;
    END
  END Address[800]
  PIN Address[801]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1335.560 4.000 1336.160 ;
    END
  END Address[801]
  PIN Address[802]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1339.640 4.000 1340.240 ;
    END
  END Address[802]
  PIN Address[803]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1343.720 4.000 1344.320 ;
    END
  END Address[803]
  PIN Address[804]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1347.800 4.000 1348.400 ;
    END
  END Address[804]
  PIN Address[805]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1351.880 4.000 1352.480 ;
    END
  END Address[805]
  PIN Address[806]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1355.960 4.000 1356.560 ;
    END
  END Address[806]
  PIN Address[807]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1360.040 4.000 1360.640 ;
    END
  END Address[807]
  PIN Address[808]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1364.120 4.000 1364.720 ;
    END
  END Address[808]
  PIN Address[809]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1368.200 4.000 1368.800 ;
    END
  END Address[809]
  PIN Address[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 482.840 800.000 483.440 ;
    END
  END Address[80]
  PIN Address[810]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1372.280 4.000 1372.880 ;
    END
  END Address[810]
  PIN Address[811]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1376.360 4.000 1376.960 ;
    END
  END Address[811]
  PIN Address[812]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1380.440 4.000 1381.040 ;
    END
  END Address[812]
  PIN Address[813]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1384.520 4.000 1385.120 ;
    END
  END Address[813]
  PIN Address[814]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1388.600 4.000 1389.200 ;
    END
  END Address[814]
  PIN Address[815]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1392.680 4.000 1393.280 ;
    END
  END Address[815]
  PIN Address[816]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1396.760 4.000 1397.360 ;
    END
  END Address[816]
  PIN Address[817]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1400.840 4.000 1401.440 ;
    END
  END Address[817]
  PIN Address[818]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1404.920 4.000 1405.520 ;
    END
  END Address[818]
  PIN Address[819]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1409.000 4.000 1409.600 ;
    END
  END Address[819]
  PIN Address[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 486.920 800.000 487.520 ;
    END
  END Address[81]
  PIN Address[820]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1413.080 4.000 1413.680 ;
    END
  END Address[820]
  PIN Address[821]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1417.160 4.000 1417.760 ;
    END
  END Address[821]
  PIN Address[822]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1421.240 4.000 1421.840 ;
    END
  END Address[822]
  PIN Address[823]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1425.320 4.000 1425.920 ;
    END
  END Address[823]
  PIN Address[824]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1429.400 4.000 1430.000 ;
    END
  END Address[824]
  PIN Address[825]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1433.480 4.000 1434.080 ;
    END
  END Address[825]
  PIN Address[826]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1437.560 4.000 1438.160 ;
    END
  END Address[826]
  PIN Address[827]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1441.640 4.000 1442.240 ;
    END
  END Address[827]
  PIN Address[828]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1445.720 4.000 1446.320 ;
    END
  END Address[828]
  PIN Address[829]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1449.800 4.000 1450.400 ;
    END
  END Address[829]
  PIN Address[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 491.000 800.000 491.600 ;
    END
  END Address[82]
  PIN Address[830]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1453.880 4.000 1454.480 ;
    END
  END Address[830]
  PIN Address[831]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1457.960 4.000 1458.560 ;
    END
  END Address[831]
  PIN Address[832]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1462.040 4.000 1462.640 ;
    END
  END Address[832]
  PIN Address[833]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1466.120 4.000 1466.720 ;
    END
  END Address[833]
  PIN Address[834]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1470.200 4.000 1470.800 ;
    END
  END Address[834]
  PIN Address[835]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1474.280 4.000 1474.880 ;
    END
  END Address[835]
  PIN Address[836]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1478.360 4.000 1478.960 ;
    END
  END Address[836]
  PIN Address[837]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1482.440 4.000 1483.040 ;
    END
  END Address[837]
  PIN Address[838]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1486.520 4.000 1487.120 ;
    END
  END Address[838]
  PIN Address[839]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1490.600 4.000 1491.200 ;
    END
  END Address[839]
  PIN Address[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 495.080 800.000 495.680 ;
    END
  END Address[83]
  PIN Address[840]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1494.680 4.000 1495.280 ;
    END
  END Address[840]
  PIN Address[841]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1498.760 4.000 1499.360 ;
    END
  END Address[841]
  PIN Address[842]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1502.840 4.000 1503.440 ;
    END
  END Address[842]
  PIN Address[843]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1506.920 4.000 1507.520 ;
    END
  END Address[843]
  PIN Address[844]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1511.000 4.000 1511.600 ;
    END
  END Address[844]
  PIN Address[845]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1515.080 4.000 1515.680 ;
    END
  END Address[845]
  PIN Address[846]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1519.160 4.000 1519.760 ;
    END
  END Address[846]
  PIN Address[847]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1523.240 4.000 1523.840 ;
    END
  END Address[847]
  PIN Address[848]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1527.320 4.000 1527.920 ;
    END
  END Address[848]
  PIN Address[849]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1531.400 4.000 1532.000 ;
    END
  END Address[849]
  PIN Address[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 499.160 800.000 499.760 ;
    END
  END Address[84]
  PIN Address[850]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1535.480 4.000 1536.080 ;
    END
  END Address[850]
  PIN Address[851]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1539.560 4.000 1540.160 ;
    END
  END Address[851]
  PIN Address[852]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1543.640 4.000 1544.240 ;
    END
  END Address[852]
  PIN Address[853]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1547.720 4.000 1548.320 ;
    END
  END Address[853]
  PIN Address[854]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1551.800 4.000 1552.400 ;
    END
  END Address[854]
  PIN Address[855]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1555.880 4.000 1556.480 ;
    END
  END Address[855]
  PIN Address[856]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1559.960 4.000 1560.560 ;
    END
  END Address[856]
  PIN Address[857]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1564.040 4.000 1564.640 ;
    END
  END Address[857]
  PIN Address[858]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1568.120 4.000 1568.720 ;
    END
  END Address[858]
  PIN Address[859]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1572.200 4.000 1572.800 ;
    END
  END Address[859]
  PIN Address[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 503.240 800.000 503.840 ;
    END
  END Address[85]
  PIN Address[860]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1576.280 4.000 1576.880 ;
    END
  END Address[860]
  PIN Address[861]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1580.360 4.000 1580.960 ;
    END
  END Address[861]
  PIN Address[862]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1584.440 4.000 1585.040 ;
    END
  END Address[862]
  PIN Address[863]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1588.520 4.000 1589.120 ;
    END
  END Address[863]
  PIN Address[864]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1592.600 4.000 1593.200 ;
    END
  END Address[864]
  PIN Address[865]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1596.680 4.000 1597.280 ;
    END
  END Address[865]
  PIN Address[866]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1600.760 4.000 1601.360 ;
    END
  END Address[866]
  PIN Address[867]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1604.840 4.000 1605.440 ;
    END
  END Address[867]
  PIN Address[868]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1608.920 4.000 1609.520 ;
    END
  END Address[868]
  PIN Address[869]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1613.000 4.000 1613.600 ;
    END
  END Address[869]
  PIN Address[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 507.320 800.000 507.920 ;
    END
  END Address[86]
  PIN Address[870]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1617.080 4.000 1617.680 ;
    END
  END Address[870]
  PIN Address[871]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1621.160 4.000 1621.760 ;
    END
  END Address[871]
  PIN Address[872]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1625.240 4.000 1625.840 ;
    END
  END Address[872]
  PIN Address[873]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1629.320 4.000 1629.920 ;
    END
  END Address[873]
  PIN Address[874]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1633.400 4.000 1634.000 ;
    END
  END Address[874]
  PIN Address[875]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1637.480 4.000 1638.080 ;
    END
  END Address[875]
  PIN Address[876]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1641.560 4.000 1642.160 ;
    END
  END Address[876]
  PIN Address[877]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1645.640 4.000 1646.240 ;
    END
  END Address[877]
  PIN Address[878]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1649.720 4.000 1650.320 ;
    END
  END Address[878]
  PIN Address[879]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1653.800 4.000 1654.400 ;
    END
  END Address[879]
  PIN Address[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 511.400 800.000 512.000 ;
    END
  END Address[87]
  PIN Address[880]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1657.880 4.000 1658.480 ;
    END
  END Address[880]
  PIN Address[881]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1661.960 4.000 1662.560 ;
    END
  END Address[881]
  PIN Address[882]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1666.040 4.000 1666.640 ;
    END
  END Address[882]
  PIN Address[883]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1670.120 4.000 1670.720 ;
    END
  END Address[883]
  PIN Address[884]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1674.200 4.000 1674.800 ;
    END
  END Address[884]
  PIN Address[885]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1678.280 4.000 1678.880 ;
    END
  END Address[885]
  PIN Address[886]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1682.360 4.000 1682.960 ;
    END
  END Address[886]
  PIN Address[887]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1686.440 4.000 1687.040 ;
    END
  END Address[887]
  PIN Address[888]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1690.520 4.000 1691.120 ;
    END
  END Address[888]
  PIN Address[889]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1694.600 4.000 1695.200 ;
    END
  END Address[889]
  PIN Address[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 515.480 800.000 516.080 ;
    END
  END Address[88]
  PIN Address[890]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1698.680 4.000 1699.280 ;
    END
  END Address[890]
  PIN Address[891]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1702.760 4.000 1703.360 ;
    END
  END Address[891]
  PIN Address[892]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1706.840 4.000 1707.440 ;
    END
  END Address[892]
  PIN Address[893]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1710.920 4.000 1711.520 ;
    END
  END Address[893]
  PIN Address[894]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1715.000 4.000 1715.600 ;
    END
  END Address[894]
  PIN Address[895]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1719.080 4.000 1719.680 ;
    END
  END Address[895]
  PIN Address[896]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1723.160 4.000 1723.760 ;
    END
  END Address[896]
  PIN Address[897]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1727.240 4.000 1727.840 ;
    END
  END Address[897]
  PIN Address[898]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1731.320 4.000 1731.920 ;
    END
  END Address[898]
  PIN Address[899]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1735.400 4.000 1736.000 ;
    END
  END Address[899]
  PIN Address[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 519.560 800.000 520.160 ;
    END
  END Address[89]
  PIN Address[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 189.080 800.000 189.680 ;
    END
  END Address[8]
  PIN Address[900]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1739.480 4.000 1740.080 ;
    END
  END Address[900]
  PIN Address[901]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1743.560 4.000 1744.160 ;
    END
  END Address[901]
  PIN Address[902]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1747.640 4.000 1748.240 ;
    END
  END Address[902]
  PIN Address[903]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1751.720 4.000 1752.320 ;
    END
  END Address[903]
  PIN Address[904]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1755.800 4.000 1756.400 ;
    END
  END Address[904]
  PIN Address[905]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1759.880 4.000 1760.480 ;
    END
  END Address[905]
  PIN Address[906]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1763.960 4.000 1764.560 ;
    END
  END Address[906]
  PIN Address[907]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1768.040 4.000 1768.640 ;
    END
  END Address[907]
  PIN Address[908]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1772.120 4.000 1772.720 ;
    END
  END Address[908]
  PIN Address[909]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1776.200 4.000 1776.800 ;
    END
  END Address[909]
  PIN Address[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 523.640 800.000 524.240 ;
    END
  END Address[90]
  PIN Address[910]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1780.280 4.000 1780.880 ;
    END
  END Address[910]
  PIN Address[911]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1784.360 4.000 1784.960 ;
    END
  END Address[911]
  PIN Address[912]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1788.440 4.000 1789.040 ;
    END
  END Address[912]
  PIN Address[913]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1792.520 4.000 1793.120 ;
    END
  END Address[913]
  PIN Address[914]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1796.600 4.000 1797.200 ;
    END
  END Address[914]
  PIN Address[915]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1800.680 4.000 1801.280 ;
    END
  END Address[915]
  PIN Address[916]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1804.760 4.000 1805.360 ;
    END
  END Address[916]
  PIN Address[917]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1808.840 4.000 1809.440 ;
    END
  END Address[917]
  PIN Address[918]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1812.920 4.000 1813.520 ;
    END
  END Address[918]
  PIN Address[919]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1817.000 4.000 1817.600 ;
    END
  END Address[919]
  PIN Address[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 527.720 800.000 528.320 ;
    END
  END Address[91]
  PIN Address[920]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1821.080 4.000 1821.680 ;
    END
  END Address[920]
  PIN Address[921]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1825.160 4.000 1825.760 ;
    END
  END Address[921]
  PIN Address[922]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1829.240 4.000 1829.840 ;
    END
  END Address[922]
  PIN Address[923]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1833.320 4.000 1833.920 ;
    END
  END Address[923]
  PIN Address[924]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1837.400 4.000 1838.000 ;
    END
  END Address[924]
  PIN Address[925]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1841.480 4.000 1842.080 ;
    END
  END Address[925]
  PIN Address[926]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1845.560 4.000 1846.160 ;
    END
  END Address[926]
  PIN Address[927]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1849.640 4.000 1850.240 ;
    END
  END Address[927]
  PIN Address[928]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1853.720 4.000 1854.320 ;
    END
  END Address[928]
  PIN Address[929]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1857.800 4.000 1858.400 ;
    END
  END Address[929]
  PIN Address[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 531.800 800.000 532.400 ;
    END
  END Address[92]
  PIN Address[930]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1861.880 4.000 1862.480 ;
    END
  END Address[930]
  PIN Address[931]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1865.960 4.000 1866.560 ;
    END
  END Address[931]
  PIN Address[932]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1870.040 4.000 1870.640 ;
    END
  END Address[932]
  PIN Address[933]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1874.120 4.000 1874.720 ;
    END
  END Address[933]
  PIN Address[934]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1878.200 4.000 1878.800 ;
    END
  END Address[934]
  PIN Address[935]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1882.280 4.000 1882.880 ;
    END
  END Address[935]
  PIN Address[936]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1886.360 4.000 1886.960 ;
    END
  END Address[936]
  PIN Address[937]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1890.440 4.000 1891.040 ;
    END
  END Address[937]
  PIN Address[938]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1894.520 4.000 1895.120 ;
    END
  END Address[938]
  PIN Address[939]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1898.600 4.000 1899.200 ;
    END
  END Address[939]
  PIN Address[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 535.880 800.000 536.480 ;
    END
  END Address[93]
  PIN Address[940]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1902.680 4.000 1903.280 ;
    END
  END Address[940]
  PIN Address[941]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1906.760 4.000 1907.360 ;
    END
  END Address[941]
  PIN Address[942]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1910.840 4.000 1911.440 ;
    END
  END Address[942]
  PIN Address[943]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1914.920 4.000 1915.520 ;
    END
  END Address[943]
  PIN Address[944]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1919.000 4.000 1919.600 ;
    END
  END Address[944]
  PIN Address[945]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1923.080 4.000 1923.680 ;
    END
  END Address[945]
  PIN Address[946]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1927.160 4.000 1927.760 ;
    END
  END Address[946]
  PIN Address[947]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1931.240 4.000 1931.840 ;
    END
  END Address[947]
  PIN Address[948]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1935.320 4.000 1935.920 ;
    END
  END Address[948]
  PIN Address[949]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1939.400 4.000 1940.000 ;
    END
  END Address[949]
  PIN Address[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 539.960 800.000 540.560 ;
    END
  END Address[94]
  PIN Address[950]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1943.480 4.000 1944.080 ;
    END
  END Address[950]
  PIN Address[951]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1947.560 4.000 1948.160 ;
    END
  END Address[951]
  PIN Address[952]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1951.640 4.000 1952.240 ;
    END
  END Address[952]
  PIN Address[953]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1955.720 4.000 1956.320 ;
    END
  END Address[953]
  PIN Address[954]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1959.800 4.000 1960.400 ;
    END
  END Address[954]
  PIN Address[955]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1963.880 4.000 1964.480 ;
    END
  END Address[955]
  PIN Address[956]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1967.960 4.000 1968.560 ;
    END
  END Address[956]
  PIN Address[957]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1972.040 4.000 1972.640 ;
    END
  END Address[957]
  PIN Address[958]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1976.120 4.000 1976.720 ;
    END
  END Address[958]
  PIN Address[959]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1980.200 4.000 1980.800 ;
    END
  END Address[959]
  PIN Address[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 544.040 800.000 544.640 ;
    END
  END Address[95]
  PIN Address[960]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1984.280 4.000 1984.880 ;
    END
  END Address[960]
  PIN Address[961]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1988.360 4.000 1988.960 ;
    END
  END Address[961]
  PIN Address[962]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1992.440 4.000 1993.040 ;
    END
  END Address[962]
  PIN Address[963]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1996.520 4.000 1997.120 ;
    END
  END Address[963]
  PIN Address[964]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2000.600 4.000 2001.200 ;
    END
  END Address[964]
  PIN Address[965]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2004.680 4.000 2005.280 ;
    END
  END Address[965]
  PIN Address[966]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2008.760 4.000 2009.360 ;
    END
  END Address[966]
  PIN Address[967]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2012.840 4.000 2013.440 ;
    END
  END Address[967]
  PIN Address[968]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2016.920 4.000 2017.520 ;
    END
  END Address[968]
  PIN Address[969]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2021.000 4.000 2021.600 ;
    END
  END Address[969]
  PIN Address[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 548.120 800.000 548.720 ;
    END
  END Address[96]
  PIN Address[970]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2025.080 4.000 2025.680 ;
    END
  END Address[970]
  PIN Address[971]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2029.160 4.000 2029.760 ;
    END
  END Address[971]
  PIN Address[972]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2033.240 4.000 2033.840 ;
    END
  END Address[972]
  PIN Address[973]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2037.320 4.000 2037.920 ;
    END
  END Address[973]
  PIN Address[974]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2041.400 4.000 2042.000 ;
    END
  END Address[974]
  PIN Address[975]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2045.480 4.000 2046.080 ;
    END
  END Address[975]
  PIN Address[976]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2049.560 4.000 2050.160 ;
    END
  END Address[976]
  PIN Address[977]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2053.640 4.000 2054.240 ;
    END
  END Address[977]
  PIN Address[978]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2057.720 4.000 2058.320 ;
    END
  END Address[978]
  PIN Address[979]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2061.800 4.000 2062.400 ;
    END
  END Address[979]
  PIN Address[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 552.200 800.000 552.800 ;
    END
  END Address[97]
  PIN Address[980]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2065.880 4.000 2066.480 ;
    END
  END Address[980]
  PIN Address[981]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2069.960 4.000 2070.560 ;
    END
  END Address[981]
  PIN Address[982]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2074.040 4.000 2074.640 ;
    END
  END Address[982]
  PIN Address[983]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2078.120 4.000 2078.720 ;
    END
  END Address[983]
  PIN Address[984]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2082.200 4.000 2082.800 ;
    END
  END Address[984]
  PIN Address[985]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2086.280 4.000 2086.880 ;
    END
  END Address[985]
  PIN Address[986]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2090.360 4.000 2090.960 ;
    END
  END Address[986]
  PIN Address[987]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2094.440 4.000 2095.040 ;
    END
  END Address[987]
  PIN Address[988]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2098.520 4.000 2099.120 ;
    END
  END Address[988]
  PIN Address[989]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2102.600 4.000 2103.200 ;
    END
  END Address[989]
  PIN Address[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 556.280 800.000 556.880 ;
    END
  END Address[98]
  PIN Address[990]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2106.680 4.000 2107.280 ;
    END
  END Address[990]
  PIN Address[991]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2110.760 4.000 2111.360 ;
    END
  END Address[991]
  PIN Address[992]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2114.840 4.000 2115.440 ;
    END
  END Address[992]
  PIN Address[993]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2118.920 4.000 2119.520 ;
    END
  END Address[993]
  PIN Address[994]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2123.000 4.000 2123.600 ;
    END
  END Address[994]
  PIN Address[995]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2127.080 4.000 2127.680 ;
    END
  END Address[995]
  PIN Address[996]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2131.160 4.000 2131.760 ;
    END
  END Address[996]
  PIN Address[997]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2135.240 4.000 2135.840 ;
    END
  END Address[997]
  PIN Address[998]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2139.320 4.000 2139.920 ;
    END
  END Address[998]
  PIN Address[999]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2143.400 4.000 2144.000 ;
    END
  END Address[999]
  PIN Address[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 560.360 800.000 560.960 ;
    END
  END Address[99]
  PIN Address[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 796.000 193.160 800.000 193.760 ;
    END
  END Address[9]
  PIN DataIn[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 8.370 2396.000 8.650 2400.000 ;
    END
  END DataIn[0]
  PIN DataIn[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 256.770 2396.000 257.050 2400.000 ;
    END
  END DataIn[10]
  PIN DataIn[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 281.610 2396.000 281.890 2400.000 ;
    END
  END DataIn[11]
  PIN DataIn[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 306.450 2396.000 306.730 2400.000 ;
    END
  END DataIn[12]
  PIN DataIn[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 331.290 2396.000 331.570 2400.000 ;
    END
  END DataIn[13]
  PIN DataIn[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 356.130 2396.000 356.410 2400.000 ;
    END
  END DataIn[14]
  PIN DataIn[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 380.970 2396.000 381.250 2400.000 ;
    END
  END DataIn[15]
  PIN DataIn[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 405.810 2396.000 406.090 2400.000 ;
    END
  END DataIn[16]
  PIN DataIn[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 430.650 2396.000 430.930 2400.000 ;
    END
  END DataIn[17]
  PIN DataIn[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 455.490 2396.000 455.770 2400.000 ;
    END
  END DataIn[18]
  PIN DataIn[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 480.330 2396.000 480.610 2400.000 ;
    END
  END DataIn[19]
  PIN DataIn[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 33.210 2396.000 33.490 2400.000 ;
    END
  END DataIn[1]
  PIN DataIn[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 505.170 2396.000 505.450 2400.000 ;
    END
  END DataIn[20]
  PIN DataIn[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 530.010 2396.000 530.290 2400.000 ;
    END
  END DataIn[21]
  PIN DataIn[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 554.850 2396.000 555.130 2400.000 ;
    END
  END DataIn[22]
  PIN DataIn[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 579.690 2396.000 579.970 2400.000 ;
    END
  END DataIn[23]
  PIN DataIn[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 604.530 2396.000 604.810 2400.000 ;
    END
  END DataIn[24]
  PIN DataIn[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 629.370 2396.000 629.650 2400.000 ;
    END
  END DataIn[25]
  PIN DataIn[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 654.210 2396.000 654.490 2400.000 ;
    END
  END DataIn[26]
  PIN DataIn[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 679.050 2396.000 679.330 2400.000 ;
    END
  END DataIn[27]
  PIN DataIn[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 703.890 2396.000 704.170 2400.000 ;
    END
  END DataIn[28]
  PIN DataIn[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 728.730 2396.000 729.010 2400.000 ;
    END
  END DataIn[29]
  PIN DataIn[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 58.050 2396.000 58.330 2400.000 ;
    END
  END DataIn[2]
  PIN DataIn[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 753.570 2396.000 753.850 2400.000 ;
    END
  END DataIn[30]
  PIN DataIn[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 778.410 2396.000 778.690 2400.000 ;
    END
  END DataIn[31]
  PIN DataIn[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 82.890 2396.000 83.170 2400.000 ;
    END
  END DataIn[3]
  PIN DataIn[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 107.730 2396.000 108.010 2400.000 ;
    END
  END DataIn[4]
  PIN DataIn[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 132.570 2396.000 132.850 2400.000 ;
    END
  END DataIn[5]
  PIN DataIn[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 157.410 2396.000 157.690 2400.000 ;
    END
  END DataIn[6]
  PIN DataIn[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 182.250 2396.000 182.530 2400.000 ;
    END
  END DataIn[7]
  PIN DataIn[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 207.090 2396.000 207.370 2400.000 ;
    END
  END DataIn[8]
  PIN DataIn[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 231.930 2396.000 232.210 2400.000 ;
    END
  END DataIn[9]
  PIN DataOut[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 20.790 2396.000 21.070 2400.000 ;
    END
  END DataOut[0]
  PIN DataOut[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 269.190 2396.000 269.470 2400.000 ;
    END
  END DataOut[10]
  PIN DataOut[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 294.030 2396.000 294.310 2400.000 ;
    END
  END DataOut[11]
  PIN DataOut[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 318.870 2396.000 319.150 2400.000 ;
    END
  END DataOut[12]
  PIN DataOut[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 343.710 2396.000 343.990 2400.000 ;
    END
  END DataOut[13]
  PIN DataOut[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 368.550 2396.000 368.830 2400.000 ;
    END
  END DataOut[14]
  PIN DataOut[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 393.390 2396.000 393.670 2400.000 ;
    END
  END DataOut[15]
  PIN DataOut[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 418.230 2396.000 418.510 2400.000 ;
    END
  END DataOut[16]
  PIN DataOut[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 443.070 2396.000 443.350 2400.000 ;
    END
  END DataOut[17]
  PIN DataOut[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 467.910 2396.000 468.190 2400.000 ;
    END
  END DataOut[18]
  PIN DataOut[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 492.750 2396.000 493.030 2400.000 ;
    END
  END DataOut[19]
  PIN DataOut[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 45.630 2396.000 45.910 2400.000 ;
    END
  END DataOut[1]
  PIN DataOut[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 517.590 2396.000 517.870 2400.000 ;
    END
  END DataOut[20]
  PIN DataOut[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 542.430 2396.000 542.710 2400.000 ;
    END
  END DataOut[21]
  PIN DataOut[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 567.270 2396.000 567.550 2400.000 ;
    END
  END DataOut[22]
  PIN DataOut[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 592.110 2396.000 592.390 2400.000 ;
    END
  END DataOut[23]
  PIN DataOut[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 616.950 2396.000 617.230 2400.000 ;
    END
  END DataOut[24]
  PIN DataOut[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 641.790 2396.000 642.070 2400.000 ;
    END
  END DataOut[25]
  PIN DataOut[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 666.630 2396.000 666.910 2400.000 ;
    END
  END DataOut[26]
  PIN DataOut[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 691.470 2396.000 691.750 2400.000 ;
    END
  END DataOut[27]
  PIN DataOut[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 716.310 2396.000 716.590 2400.000 ;
    END
  END DataOut[28]
  PIN DataOut[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 741.150 2396.000 741.430 2400.000 ;
    END
  END DataOut[29]
  PIN DataOut[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 70.470 2396.000 70.750 2400.000 ;
    END
  END DataOut[2]
  PIN DataOut[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 765.990 2396.000 766.270 2400.000 ;
    END
  END DataOut[30]
  PIN DataOut[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 790.830 2396.000 791.110 2400.000 ;
    END
  END DataOut[31]
  PIN DataOut[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 95.310 2396.000 95.590 2400.000 ;
    END
  END DataOut[3]
  PIN DataOut[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 120.150 2396.000 120.430 2400.000 ;
    END
  END DataOut[4]
  PIN DataOut[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 144.990 2396.000 145.270 2400.000 ;
    END
  END DataOut[5]
  PIN DataOut[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 169.830 2396.000 170.110 2400.000 ;
    END
  END DataOut[6]
  PIN DataOut[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 194.670 2396.000 194.950 2400.000 ;
    END
  END DataOut[7]
  PIN DataOut[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 219.510 2396.000 219.790 2400.000 ;
    END
  END DataOut[8]
  PIN DataOut[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 244.350 2396.000 244.630 2400.000 ;
    END
  END DataOut[9]
  PIN PRE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 133.490 0.000 133.770 4.000 ;
    END
  END PRE
  PIN ReadEn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 399.830 0.000 400.110 4.000 ;
    END
  END ReadEn
  PIN WriteEn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 666.170 0.000 666.450 4.000 ;
    END
  END WriteEn
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 2388.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 2388.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 2388.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 2388.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 2388.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 2388.400 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 2388.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 2388.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 2388.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 2388.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 2388.400 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 795.195 2388.245 ;
      LAYER met1 ;
        RECT 1.910 10.640 798.490 2388.400 ;
      LAYER met2 ;
        RECT 1.930 2395.720 8.090 2396.730 ;
        RECT 8.930 2395.720 20.510 2396.730 ;
        RECT 21.350 2395.720 32.930 2396.730 ;
        RECT 33.770 2395.720 45.350 2396.730 ;
        RECT 46.190 2395.720 57.770 2396.730 ;
        RECT 58.610 2395.720 70.190 2396.730 ;
        RECT 71.030 2395.720 82.610 2396.730 ;
        RECT 83.450 2395.720 95.030 2396.730 ;
        RECT 95.870 2395.720 107.450 2396.730 ;
        RECT 108.290 2395.720 119.870 2396.730 ;
        RECT 120.710 2395.720 132.290 2396.730 ;
        RECT 133.130 2395.720 144.710 2396.730 ;
        RECT 145.550 2395.720 157.130 2396.730 ;
        RECT 157.970 2395.720 169.550 2396.730 ;
        RECT 170.390 2395.720 181.970 2396.730 ;
        RECT 182.810 2395.720 194.390 2396.730 ;
        RECT 195.230 2395.720 206.810 2396.730 ;
        RECT 207.650 2395.720 219.230 2396.730 ;
        RECT 220.070 2395.720 231.650 2396.730 ;
        RECT 232.490 2395.720 244.070 2396.730 ;
        RECT 244.910 2395.720 256.490 2396.730 ;
        RECT 257.330 2395.720 268.910 2396.730 ;
        RECT 269.750 2395.720 281.330 2396.730 ;
        RECT 282.170 2395.720 293.750 2396.730 ;
        RECT 294.590 2395.720 306.170 2396.730 ;
        RECT 307.010 2395.720 318.590 2396.730 ;
        RECT 319.430 2395.720 331.010 2396.730 ;
        RECT 331.850 2395.720 343.430 2396.730 ;
        RECT 344.270 2395.720 355.850 2396.730 ;
        RECT 356.690 2395.720 368.270 2396.730 ;
        RECT 369.110 2395.720 380.690 2396.730 ;
        RECT 381.530 2395.720 393.110 2396.730 ;
        RECT 393.950 2395.720 405.530 2396.730 ;
        RECT 406.370 2395.720 417.950 2396.730 ;
        RECT 418.790 2395.720 430.370 2396.730 ;
        RECT 431.210 2395.720 442.790 2396.730 ;
        RECT 443.630 2395.720 455.210 2396.730 ;
        RECT 456.050 2395.720 467.630 2396.730 ;
        RECT 468.470 2395.720 480.050 2396.730 ;
        RECT 480.890 2395.720 492.470 2396.730 ;
        RECT 493.310 2395.720 504.890 2396.730 ;
        RECT 505.730 2395.720 517.310 2396.730 ;
        RECT 518.150 2395.720 529.730 2396.730 ;
        RECT 530.570 2395.720 542.150 2396.730 ;
        RECT 542.990 2395.720 554.570 2396.730 ;
        RECT 555.410 2395.720 566.990 2396.730 ;
        RECT 567.830 2395.720 579.410 2396.730 ;
        RECT 580.250 2395.720 591.830 2396.730 ;
        RECT 592.670 2395.720 604.250 2396.730 ;
        RECT 605.090 2395.720 616.670 2396.730 ;
        RECT 617.510 2395.720 629.090 2396.730 ;
        RECT 629.930 2395.720 641.510 2396.730 ;
        RECT 642.350 2395.720 653.930 2396.730 ;
        RECT 654.770 2395.720 666.350 2396.730 ;
        RECT 667.190 2395.720 678.770 2396.730 ;
        RECT 679.610 2395.720 691.190 2396.730 ;
        RECT 692.030 2395.720 703.610 2396.730 ;
        RECT 704.450 2395.720 716.030 2396.730 ;
        RECT 716.870 2395.720 728.450 2396.730 ;
        RECT 729.290 2395.720 740.870 2396.730 ;
        RECT 741.710 2395.720 753.290 2396.730 ;
        RECT 754.130 2395.720 765.710 2396.730 ;
        RECT 766.550 2395.720 778.130 2396.730 ;
        RECT 778.970 2395.720 790.550 2396.730 ;
        RECT 791.390 2395.720 798.470 2396.730 ;
        RECT 1.930 4.280 798.470 2395.720 ;
        RECT 1.930 4.000 133.210 4.280 ;
        RECT 134.050 4.000 399.550 4.280 ;
        RECT 400.390 4.000 665.890 4.280 ;
        RECT 666.730 4.000 798.470 4.280 ;
      LAYER met3 ;
        RECT 1.905 2242.320 798.495 2388.325 ;
        RECT 4.400 2240.920 795.600 2242.320 ;
        RECT 1.905 2238.240 798.495 2240.920 ;
        RECT 4.400 2236.840 795.600 2238.240 ;
        RECT 1.905 2234.160 798.495 2236.840 ;
        RECT 4.400 2232.760 795.600 2234.160 ;
        RECT 1.905 2230.080 798.495 2232.760 ;
        RECT 4.400 2228.680 795.600 2230.080 ;
        RECT 1.905 2226.000 798.495 2228.680 ;
        RECT 4.400 2224.600 795.600 2226.000 ;
        RECT 1.905 2221.920 798.495 2224.600 ;
        RECT 4.400 2220.520 795.600 2221.920 ;
        RECT 1.905 2217.840 798.495 2220.520 ;
        RECT 4.400 2216.440 795.600 2217.840 ;
        RECT 1.905 2213.760 798.495 2216.440 ;
        RECT 4.400 2212.360 795.600 2213.760 ;
        RECT 1.905 2209.680 798.495 2212.360 ;
        RECT 4.400 2208.280 795.600 2209.680 ;
        RECT 1.905 2205.600 798.495 2208.280 ;
        RECT 4.400 2204.200 795.600 2205.600 ;
        RECT 1.905 2201.520 798.495 2204.200 ;
        RECT 4.400 2200.120 795.600 2201.520 ;
        RECT 1.905 2197.440 798.495 2200.120 ;
        RECT 4.400 2196.040 795.600 2197.440 ;
        RECT 1.905 2193.360 798.495 2196.040 ;
        RECT 4.400 2191.960 795.600 2193.360 ;
        RECT 1.905 2189.280 798.495 2191.960 ;
        RECT 4.400 2187.880 795.600 2189.280 ;
        RECT 1.905 2185.200 798.495 2187.880 ;
        RECT 4.400 2183.800 795.600 2185.200 ;
        RECT 1.905 2181.120 798.495 2183.800 ;
        RECT 4.400 2179.720 795.600 2181.120 ;
        RECT 1.905 2177.040 798.495 2179.720 ;
        RECT 4.400 2175.640 795.600 2177.040 ;
        RECT 1.905 2172.960 798.495 2175.640 ;
        RECT 4.400 2171.560 795.600 2172.960 ;
        RECT 1.905 2168.880 798.495 2171.560 ;
        RECT 4.400 2167.480 795.600 2168.880 ;
        RECT 1.905 2164.800 798.495 2167.480 ;
        RECT 4.400 2163.400 795.600 2164.800 ;
        RECT 1.905 2160.720 798.495 2163.400 ;
        RECT 4.400 2159.320 795.600 2160.720 ;
        RECT 1.905 2156.640 798.495 2159.320 ;
        RECT 4.400 2155.240 795.600 2156.640 ;
        RECT 1.905 2152.560 798.495 2155.240 ;
        RECT 4.400 2151.160 795.600 2152.560 ;
        RECT 1.905 2148.480 798.495 2151.160 ;
        RECT 4.400 2147.080 795.600 2148.480 ;
        RECT 1.905 2144.400 798.495 2147.080 ;
        RECT 4.400 2143.000 795.600 2144.400 ;
        RECT 1.905 2140.320 798.495 2143.000 ;
        RECT 4.400 2138.920 795.600 2140.320 ;
        RECT 1.905 2136.240 798.495 2138.920 ;
        RECT 4.400 2134.840 795.600 2136.240 ;
        RECT 1.905 2132.160 798.495 2134.840 ;
        RECT 4.400 2130.760 795.600 2132.160 ;
        RECT 1.905 2128.080 798.495 2130.760 ;
        RECT 4.400 2126.680 795.600 2128.080 ;
        RECT 1.905 2124.000 798.495 2126.680 ;
        RECT 4.400 2122.600 795.600 2124.000 ;
        RECT 1.905 2119.920 798.495 2122.600 ;
        RECT 4.400 2118.520 795.600 2119.920 ;
        RECT 1.905 2115.840 798.495 2118.520 ;
        RECT 4.400 2114.440 795.600 2115.840 ;
        RECT 1.905 2111.760 798.495 2114.440 ;
        RECT 4.400 2110.360 795.600 2111.760 ;
        RECT 1.905 2107.680 798.495 2110.360 ;
        RECT 4.400 2106.280 795.600 2107.680 ;
        RECT 1.905 2103.600 798.495 2106.280 ;
        RECT 4.400 2102.200 795.600 2103.600 ;
        RECT 1.905 2099.520 798.495 2102.200 ;
        RECT 4.400 2098.120 795.600 2099.520 ;
        RECT 1.905 2095.440 798.495 2098.120 ;
        RECT 4.400 2094.040 795.600 2095.440 ;
        RECT 1.905 2091.360 798.495 2094.040 ;
        RECT 4.400 2089.960 795.600 2091.360 ;
        RECT 1.905 2087.280 798.495 2089.960 ;
        RECT 4.400 2085.880 795.600 2087.280 ;
        RECT 1.905 2083.200 798.495 2085.880 ;
        RECT 4.400 2081.800 795.600 2083.200 ;
        RECT 1.905 2079.120 798.495 2081.800 ;
        RECT 4.400 2077.720 795.600 2079.120 ;
        RECT 1.905 2075.040 798.495 2077.720 ;
        RECT 4.400 2073.640 795.600 2075.040 ;
        RECT 1.905 2070.960 798.495 2073.640 ;
        RECT 4.400 2069.560 795.600 2070.960 ;
        RECT 1.905 2066.880 798.495 2069.560 ;
        RECT 4.400 2065.480 795.600 2066.880 ;
        RECT 1.905 2062.800 798.495 2065.480 ;
        RECT 4.400 2061.400 795.600 2062.800 ;
        RECT 1.905 2058.720 798.495 2061.400 ;
        RECT 4.400 2057.320 795.600 2058.720 ;
        RECT 1.905 2054.640 798.495 2057.320 ;
        RECT 4.400 2053.240 795.600 2054.640 ;
        RECT 1.905 2050.560 798.495 2053.240 ;
        RECT 4.400 2049.160 795.600 2050.560 ;
        RECT 1.905 2046.480 798.495 2049.160 ;
        RECT 4.400 2045.080 795.600 2046.480 ;
        RECT 1.905 2042.400 798.495 2045.080 ;
        RECT 4.400 2041.000 795.600 2042.400 ;
        RECT 1.905 2038.320 798.495 2041.000 ;
        RECT 4.400 2036.920 795.600 2038.320 ;
        RECT 1.905 2034.240 798.495 2036.920 ;
        RECT 4.400 2032.840 795.600 2034.240 ;
        RECT 1.905 2030.160 798.495 2032.840 ;
        RECT 4.400 2028.760 795.600 2030.160 ;
        RECT 1.905 2026.080 798.495 2028.760 ;
        RECT 4.400 2024.680 795.600 2026.080 ;
        RECT 1.905 2022.000 798.495 2024.680 ;
        RECT 4.400 2020.600 795.600 2022.000 ;
        RECT 1.905 2017.920 798.495 2020.600 ;
        RECT 4.400 2016.520 795.600 2017.920 ;
        RECT 1.905 2013.840 798.495 2016.520 ;
        RECT 4.400 2012.440 795.600 2013.840 ;
        RECT 1.905 2009.760 798.495 2012.440 ;
        RECT 4.400 2008.360 795.600 2009.760 ;
        RECT 1.905 2005.680 798.495 2008.360 ;
        RECT 4.400 2004.280 795.600 2005.680 ;
        RECT 1.905 2001.600 798.495 2004.280 ;
        RECT 4.400 2000.200 795.600 2001.600 ;
        RECT 1.905 1997.520 798.495 2000.200 ;
        RECT 4.400 1996.120 795.600 1997.520 ;
        RECT 1.905 1993.440 798.495 1996.120 ;
        RECT 4.400 1992.040 795.600 1993.440 ;
        RECT 1.905 1989.360 798.495 1992.040 ;
        RECT 4.400 1987.960 795.600 1989.360 ;
        RECT 1.905 1985.280 798.495 1987.960 ;
        RECT 4.400 1983.880 795.600 1985.280 ;
        RECT 1.905 1981.200 798.495 1983.880 ;
        RECT 4.400 1979.800 795.600 1981.200 ;
        RECT 1.905 1977.120 798.495 1979.800 ;
        RECT 4.400 1975.720 795.600 1977.120 ;
        RECT 1.905 1973.040 798.495 1975.720 ;
        RECT 4.400 1971.640 795.600 1973.040 ;
        RECT 1.905 1968.960 798.495 1971.640 ;
        RECT 4.400 1967.560 795.600 1968.960 ;
        RECT 1.905 1964.880 798.495 1967.560 ;
        RECT 4.400 1963.480 795.600 1964.880 ;
        RECT 1.905 1960.800 798.495 1963.480 ;
        RECT 4.400 1959.400 795.600 1960.800 ;
        RECT 1.905 1956.720 798.495 1959.400 ;
        RECT 4.400 1955.320 795.600 1956.720 ;
        RECT 1.905 1952.640 798.495 1955.320 ;
        RECT 4.400 1951.240 795.600 1952.640 ;
        RECT 1.905 1948.560 798.495 1951.240 ;
        RECT 4.400 1947.160 795.600 1948.560 ;
        RECT 1.905 1944.480 798.495 1947.160 ;
        RECT 4.400 1943.080 795.600 1944.480 ;
        RECT 1.905 1940.400 798.495 1943.080 ;
        RECT 4.400 1939.000 795.600 1940.400 ;
        RECT 1.905 1936.320 798.495 1939.000 ;
        RECT 4.400 1934.920 795.600 1936.320 ;
        RECT 1.905 1932.240 798.495 1934.920 ;
        RECT 4.400 1930.840 795.600 1932.240 ;
        RECT 1.905 1928.160 798.495 1930.840 ;
        RECT 4.400 1926.760 795.600 1928.160 ;
        RECT 1.905 1924.080 798.495 1926.760 ;
        RECT 4.400 1922.680 795.600 1924.080 ;
        RECT 1.905 1920.000 798.495 1922.680 ;
        RECT 4.400 1918.600 795.600 1920.000 ;
        RECT 1.905 1915.920 798.495 1918.600 ;
        RECT 4.400 1914.520 795.600 1915.920 ;
        RECT 1.905 1911.840 798.495 1914.520 ;
        RECT 4.400 1910.440 795.600 1911.840 ;
        RECT 1.905 1907.760 798.495 1910.440 ;
        RECT 4.400 1906.360 795.600 1907.760 ;
        RECT 1.905 1903.680 798.495 1906.360 ;
        RECT 4.400 1902.280 795.600 1903.680 ;
        RECT 1.905 1899.600 798.495 1902.280 ;
        RECT 4.400 1898.200 795.600 1899.600 ;
        RECT 1.905 1895.520 798.495 1898.200 ;
        RECT 4.400 1894.120 795.600 1895.520 ;
        RECT 1.905 1891.440 798.495 1894.120 ;
        RECT 4.400 1890.040 795.600 1891.440 ;
        RECT 1.905 1887.360 798.495 1890.040 ;
        RECT 4.400 1885.960 795.600 1887.360 ;
        RECT 1.905 1883.280 798.495 1885.960 ;
        RECT 4.400 1881.880 795.600 1883.280 ;
        RECT 1.905 1879.200 798.495 1881.880 ;
        RECT 4.400 1877.800 795.600 1879.200 ;
        RECT 1.905 1875.120 798.495 1877.800 ;
        RECT 4.400 1873.720 795.600 1875.120 ;
        RECT 1.905 1871.040 798.495 1873.720 ;
        RECT 4.400 1869.640 795.600 1871.040 ;
        RECT 1.905 1866.960 798.495 1869.640 ;
        RECT 4.400 1865.560 795.600 1866.960 ;
        RECT 1.905 1862.880 798.495 1865.560 ;
        RECT 4.400 1861.480 795.600 1862.880 ;
        RECT 1.905 1858.800 798.495 1861.480 ;
        RECT 4.400 1857.400 795.600 1858.800 ;
        RECT 1.905 1854.720 798.495 1857.400 ;
        RECT 4.400 1853.320 795.600 1854.720 ;
        RECT 1.905 1850.640 798.495 1853.320 ;
        RECT 4.400 1849.240 795.600 1850.640 ;
        RECT 1.905 1846.560 798.495 1849.240 ;
        RECT 4.400 1845.160 795.600 1846.560 ;
        RECT 1.905 1842.480 798.495 1845.160 ;
        RECT 4.400 1841.080 795.600 1842.480 ;
        RECT 1.905 1838.400 798.495 1841.080 ;
        RECT 4.400 1837.000 795.600 1838.400 ;
        RECT 1.905 1834.320 798.495 1837.000 ;
        RECT 4.400 1832.920 795.600 1834.320 ;
        RECT 1.905 1830.240 798.495 1832.920 ;
        RECT 4.400 1828.840 795.600 1830.240 ;
        RECT 1.905 1826.160 798.495 1828.840 ;
        RECT 4.400 1824.760 795.600 1826.160 ;
        RECT 1.905 1822.080 798.495 1824.760 ;
        RECT 4.400 1820.680 795.600 1822.080 ;
        RECT 1.905 1818.000 798.495 1820.680 ;
        RECT 4.400 1816.600 795.600 1818.000 ;
        RECT 1.905 1813.920 798.495 1816.600 ;
        RECT 4.400 1812.520 795.600 1813.920 ;
        RECT 1.905 1809.840 798.495 1812.520 ;
        RECT 4.400 1808.440 795.600 1809.840 ;
        RECT 1.905 1805.760 798.495 1808.440 ;
        RECT 4.400 1804.360 795.600 1805.760 ;
        RECT 1.905 1801.680 798.495 1804.360 ;
        RECT 4.400 1800.280 795.600 1801.680 ;
        RECT 1.905 1797.600 798.495 1800.280 ;
        RECT 4.400 1796.200 795.600 1797.600 ;
        RECT 1.905 1793.520 798.495 1796.200 ;
        RECT 4.400 1792.120 795.600 1793.520 ;
        RECT 1.905 1789.440 798.495 1792.120 ;
        RECT 4.400 1788.040 795.600 1789.440 ;
        RECT 1.905 1785.360 798.495 1788.040 ;
        RECT 4.400 1783.960 795.600 1785.360 ;
        RECT 1.905 1781.280 798.495 1783.960 ;
        RECT 4.400 1779.880 795.600 1781.280 ;
        RECT 1.905 1777.200 798.495 1779.880 ;
        RECT 4.400 1775.800 795.600 1777.200 ;
        RECT 1.905 1773.120 798.495 1775.800 ;
        RECT 4.400 1771.720 795.600 1773.120 ;
        RECT 1.905 1769.040 798.495 1771.720 ;
        RECT 4.400 1767.640 795.600 1769.040 ;
        RECT 1.905 1764.960 798.495 1767.640 ;
        RECT 4.400 1763.560 795.600 1764.960 ;
        RECT 1.905 1760.880 798.495 1763.560 ;
        RECT 4.400 1759.480 795.600 1760.880 ;
        RECT 1.905 1756.800 798.495 1759.480 ;
        RECT 4.400 1755.400 795.600 1756.800 ;
        RECT 1.905 1752.720 798.495 1755.400 ;
        RECT 4.400 1751.320 795.600 1752.720 ;
        RECT 1.905 1748.640 798.495 1751.320 ;
        RECT 4.400 1747.240 795.600 1748.640 ;
        RECT 1.905 1744.560 798.495 1747.240 ;
        RECT 4.400 1743.160 795.600 1744.560 ;
        RECT 1.905 1740.480 798.495 1743.160 ;
        RECT 4.400 1739.080 795.600 1740.480 ;
        RECT 1.905 1736.400 798.495 1739.080 ;
        RECT 4.400 1735.000 795.600 1736.400 ;
        RECT 1.905 1732.320 798.495 1735.000 ;
        RECT 4.400 1730.920 795.600 1732.320 ;
        RECT 1.905 1728.240 798.495 1730.920 ;
        RECT 4.400 1726.840 795.600 1728.240 ;
        RECT 1.905 1724.160 798.495 1726.840 ;
        RECT 4.400 1722.760 795.600 1724.160 ;
        RECT 1.905 1720.080 798.495 1722.760 ;
        RECT 4.400 1718.680 795.600 1720.080 ;
        RECT 1.905 1716.000 798.495 1718.680 ;
        RECT 4.400 1714.600 795.600 1716.000 ;
        RECT 1.905 1711.920 798.495 1714.600 ;
        RECT 4.400 1710.520 795.600 1711.920 ;
        RECT 1.905 1707.840 798.495 1710.520 ;
        RECT 4.400 1706.440 795.600 1707.840 ;
        RECT 1.905 1703.760 798.495 1706.440 ;
        RECT 4.400 1702.360 795.600 1703.760 ;
        RECT 1.905 1699.680 798.495 1702.360 ;
        RECT 4.400 1698.280 795.600 1699.680 ;
        RECT 1.905 1695.600 798.495 1698.280 ;
        RECT 4.400 1694.200 795.600 1695.600 ;
        RECT 1.905 1691.520 798.495 1694.200 ;
        RECT 4.400 1690.120 795.600 1691.520 ;
        RECT 1.905 1687.440 798.495 1690.120 ;
        RECT 4.400 1686.040 795.600 1687.440 ;
        RECT 1.905 1683.360 798.495 1686.040 ;
        RECT 4.400 1681.960 795.600 1683.360 ;
        RECT 1.905 1679.280 798.495 1681.960 ;
        RECT 4.400 1677.880 795.600 1679.280 ;
        RECT 1.905 1675.200 798.495 1677.880 ;
        RECT 4.400 1673.800 795.600 1675.200 ;
        RECT 1.905 1671.120 798.495 1673.800 ;
        RECT 4.400 1669.720 795.600 1671.120 ;
        RECT 1.905 1667.040 798.495 1669.720 ;
        RECT 4.400 1665.640 795.600 1667.040 ;
        RECT 1.905 1662.960 798.495 1665.640 ;
        RECT 4.400 1661.560 795.600 1662.960 ;
        RECT 1.905 1658.880 798.495 1661.560 ;
        RECT 4.400 1657.480 795.600 1658.880 ;
        RECT 1.905 1654.800 798.495 1657.480 ;
        RECT 4.400 1653.400 795.600 1654.800 ;
        RECT 1.905 1650.720 798.495 1653.400 ;
        RECT 4.400 1649.320 795.600 1650.720 ;
        RECT 1.905 1646.640 798.495 1649.320 ;
        RECT 4.400 1645.240 795.600 1646.640 ;
        RECT 1.905 1642.560 798.495 1645.240 ;
        RECT 4.400 1641.160 795.600 1642.560 ;
        RECT 1.905 1638.480 798.495 1641.160 ;
        RECT 4.400 1637.080 795.600 1638.480 ;
        RECT 1.905 1634.400 798.495 1637.080 ;
        RECT 4.400 1633.000 795.600 1634.400 ;
        RECT 1.905 1630.320 798.495 1633.000 ;
        RECT 4.400 1628.920 795.600 1630.320 ;
        RECT 1.905 1626.240 798.495 1628.920 ;
        RECT 4.400 1624.840 795.600 1626.240 ;
        RECT 1.905 1622.160 798.495 1624.840 ;
        RECT 4.400 1620.760 795.600 1622.160 ;
        RECT 1.905 1618.080 798.495 1620.760 ;
        RECT 4.400 1616.680 795.600 1618.080 ;
        RECT 1.905 1614.000 798.495 1616.680 ;
        RECT 4.400 1612.600 795.600 1614.000 ;
        RECT 1.905 1609.920 798.495 1612.600 ;
        RECT 4.400 1608.520 795.600 1609.920 ;
        RECT 1.905 1605.840 798.495 1608.520 ;
        RECT 4.400 1604.440 795.600 1605.840 ;
        RECT 1.905 1601.760 798.495 1604.440 ;
        RECT 4.400 1600.360 795.600 1601.760 ;
        RECT 1.905 1597.680 798.495 1600.360 ;
        RECT 4.400 1596.280 795.600 1597.680 ;
        RECT 1.905 1593.600 798.495 1596.280 ;
        RECT 4.400 1592.200 795.600 1593.600 ;
        RECT 1.905 1589.520 798.495 1592.200 ;
        RECT 4.400 1588.120 795.600 1589.520 ;
        RECT 1.905 1585.440 798.495 1588.120 ;
        RECT 4.400 1584.040 795.600 1585.440 ;
        RECT 1.905 1581.360 798.495 1584.040 ;
        RECT 4.400 1579.960 795.600 1581.360 ;
        RECT 1.905 1577.280 798.495 1579.960 ;
        RECT 4.400 1575.880 795.600 1577.280 ;
        RECT 1.905 1573.200 798.495 1575.880 ;
        RECT 4.400 1571.800 795.600 1573.200 ;
        RECT 1.905 1569.120 798.495 1571.800 ;
        RECT 4.400 1567.720 795.600 1569.120 ;
        RECT 1.905 1565.040 798.495 1567.720 ;
        RECT 4.400 1563.640 795.600 1565.040 ;
        RECT 1.905 1560.960 798.495 1563.640 ;
        RECT 4.400 1559.560 795.600 1560.960 ;
        RECT 1.905 1556.880 798.495 1559.560 ;
        RECT 4.400 1555.480 795.600 1556.880 ;
        RECT 1.905 1552.800 798.495 1555.480 ;
        RECT 4.400 1551.400 795.600 1552.800 ;
        RECT 1.905 1548.720 798.495 1551.400 ;
        RECT 4.400 1547.320 795.600 1548.720 ;
        RECT 1.905 1544.640 798.495 1547.320 ;
        RECT 4.400 1543.240 795.600 1544.640 ;
        RECT 1.905 1540.560 798.495 1543.240 ;
        RECT 4.400 1539.160 795.600 1540.560 ;
        RECT 1.905 1536.480 798.495 1539.160 ;
        RECT 4.400 1535.080 795.600 1536.480 ;
        RECT 1.905 1532.400 798.495 1535.080 ;
        RECT 4.400 1531.000 795.600 1532.400 ;
        RECT 1.905 1528.320 798.495 1531.000 ;
        RECT 4.400 1526.920 795.600 1528.320 ;
        RECT 1.905 1524.240 798.495 1526.920 ;
        RECT 4.400 1522.840 795.600 1524.240 ;
        RECT 1.905 1520.160 798.495 1522.840 ;
        RECT 4.400 1518.760 795.600 1520.160 ;
        RECT 1.905 1516.080 798.495 1518.760 ;
        RECT 4.400 1514.680 795.600 1516.080 ;
        RECT 1.905 1512.000 798.495 1514.680 ;
        RECT 4.400 1510.600 795.600 1512.000 ;
        RECT 1.905 1507.920 798.495 1510.600 ;
        RECT 4.400 1506.520 795.600 1507.920 ;
        RECT 1.905 1503.840 798.495 1506.520 ;
        RECT 4.400 1502.440 795.600 1503.840 ;
        RECT 1.905 1499.760 798.495 1502.440 ;
        RECT 4.400 1498.360 795.600 1499.760 ;
        RECT 1.905 1495.680 798.495 1498.360 ;
        RECT 4.400 1494.280 795.600 1495.680 ;
        RECT 1.905 1491.600 798.495 1494.280 ;
        RECT 4.400 1490.200 795.600 1491.600 ;
        RECT 1.905 1487.520 798.495 1490.200 ;
        RECT 4.400 1486.120 795.600 1487.520 ;
        RECT 1.905 1483.440 798.495 1486.120 ;
        RECT 4.400 1482.040 795.600 1483.440 ;
        RECT 1.905 1479.360 798.495 1482.040 ;
        RECT 4.400 1477.960 795.600 1479.360 ;
        RECT 1.905 1475.280 798.495 1477.960 ;
        RECT 4.400 1473.880 795.600 1475.280 ;
        RECT 1.905 1471.200 798.495 1473.880 ;
        RECT 4.400 1469.800 795.600 1471.200 ;
        RECT 1.905 1467.120 798.495 1469.800 ;
        RECT 4.400 1465.720 795.600 1467.120 ;
        RECT 1.905 1463.040 798.495 1465.720 ;
        RECT 4.400 1461.640 795.600 1463.040 ;
        RECT 1.905 1458.960 798.495 1461.640 ;
        RECT 4.400 1457.560 795.600 1458.960 ;
        RECT 1.905 1454.880 798.495 1457.560 ;
        RECT 4.400 1453.480 795.600 1454.880 ;
        RECT 1.905 1450.800 798.495 1453.480 ;
        RECT 4.400 1449.400 795.600 1450.800 ;
        RECT 1.905 1446.720 798.495 1449.400 ;
        RECT 4.400 1445.320 795.600 1446.720 ;
        RECT 1.905 1442.640 798.495 1445.320 ;
        RECT 4.400 1441.240 795.600 1442.640 ;
        RECT 1.905 1438.560 798.495 1441.240 ;
        RECT 4.400 1437.160 795.600 1438.560 ;
        RECT 1.905 1434.480 798.495 1437.160 ;
        RECT 4.400 1433.080 795.600 1434.480 ;
        RECT 1.905 1430.400 798.495 1433.080 ;
        RECT 4.400 1429.000 795.600 1430.400 ;
        RECT 1.905 1426.320 798.495 1429.000 ;
        RECT 4.400 1424.920 795.600 1426.320 ;
        RECT 1.905 1422.240 798.495 1424.920 ;
        RECT 4.400 1420.840 795.600 1422.240 ;
        RECT 1.905 1418.160 798.495 1420.840 ;
        RECT 4.400 1416.760 795.600 1418.160 ;
        RECT 1.905 1414.080 798.495 1416.760 ;
        RECT 4.400 1412.680 795.600 1414.080 ;
        RECT 1.905 1410.000 798.495 1412.680 ;
        RECT 4.400 1408.600 795.600 1410.000 ;
        RECT 1.905 1405.920 798.495 1408.600 ;
        RECT 4.400 1404.520 795.600 1405.920 ;
        RECT 1.905 1401.840 798.495 1404.520 ;
        RECT 4.400 1400.440 795.600 1401.840 ;
        RECT 1.905 1397.760 798.495 1400.440 ;
        RECT 4.400 1396.360 795.600 1397.760 ;
        RECT 1.905 1393.680 798.495 1396.360 ;
        RECT 4.400 1392.280 795.600 1393.680 ;
        RECT 1.905 1389.600 798.495 1392.280 ;
        RECT 4.400 1388.200 795.600 1389.600 ;
        RECT 1.905 1385.520 798.495 1388.200 ;
        RECT 4.400 1384.120 795.600 1385.520 ;
        RECT 1.905 1381.440 798.495 1384.120 ;
        RECT 4.400 1380.040 795.600 1381.440 ;
        RECT 1.905 1377.360 798.495 1380.040 ;
        RECT 4.400 1375.960 795.600 1377.360 ;
        RECT 1.905 1373.280 798.495 1375.960 ;
        RECT 4.400 1371.880 795.600 1373.280 ;
        RECT 1.905 1369.200 798.495 1371.880 ;
        RECT 4.400 1367.800 795.600 1369.200 ;
        RECT 1.905 1365.120 798.495 1367.800 ;
        RECT 4.400 1363.720 795.600 1365.120 ;
        RECT 1.905 1361.040 798.495 1363.720 ;
        RECT 4.400 1359.640 795.600 1361.040 ;
        RECT 1.905 1356.960 798.495 1359.640 ;
        RECT 4.400 1355.560 795.600 1356.960 ;
        RECT 1.905 1352.880 798.495 1355.560 ;
        RECT 4.400 1351.480 795.600 1352.880 ;
        RECT 1.905 1348.800 798.495 1351.480 ;
        RECT 4.400 1347.400 795.600 1348.800 ;
        RECT 1.905 1344.720 798.495 1347.400 ;
        RECT 4.400 1343.320 795.600 1344.720 ;
        RECT 1.905 1340.640 798.495 1343.320 ;
        RECT 4.400 1339.240 795.600 1340.640 ;
        RECT 1.905 1336.560 798.495 1339.240 ;
        RECT 4.400 1335.160 795.600 1336.560 ;
        RECT 1.905 1332.480 798.495 1335.160 ;
        RECT 4.400 1331.080 795.600 1332.480 ;
        RECT 1.905 1328.400 798.495 1331.080 ;
        RECT 4.400 1327.000 795.600 1328.400 ;
        RECT 1.905 1324.320 798.495 1327.000 ;
        RECT 4.400 1322.920 795.600 1324.320 ;
        RECT 1.905 1320.240 798.495 1322.920 ;
        RECT 4.400 1318.840 795.600 1320.240 ;
        RECT 1.905 1316.160 798.495 1318.840 ;
        RECT 4.400 1314.760 795.600 1316.160 ;
        RECT 1.905 1312.080 798.495 1314.760 ;
        RECT 4.400 1310.680 795.600 1312.080 ;
        RECT 1.905 1308.000 798.495 1310.680 ;
        RECT 4.400 1306.600 795.600 1308.000 ;
        RECT 1.905 1303.920 798.495 1306.600 ;
        RECT 4.400 1302.520 795.600 1303.920 ;
        RECT 1.905 1299.840 798.495 1302.520 ;
        RECT 4.400 1298.440 795.600 1299.840 ;
        RECT 1.905 1295.760 798.495 1298.440 ;
        RECT 4.400 1294.360 795.600 1295.760 ;
        RECT 1.905 1291.680 798.495 1294.360 ;
        RECT 4.400 1290.280 795.600 1291.680 ;
        RECT 1.905 1287.600 798.495 1290.280 ;
        RECT 4.400 1286.200 795.600 1287.600 ;
        RECT 1.905 1283.520 798.495 1286.200 ;
        RECT 4.400 1282.120 795.600 1283.520 ;
        RECT 1.905 1279.440 798.495 1282.120 ;
        RECT 4.400 1278.040 795.600 1279.440 ;
        RECT 1.905 1275.360 798.495 1278.040 ;
        RECT 4.400 1273.960 795.600 1275.360 ;
        RECT 1.905 1271.280 798.495 1273.960 ;
        RECT 4.400 1269.880 795.600 1271.280 ;
        RECT 1.905 1267.200 798.495 1269.880 ;
        RECT 4.400 1265.800 795.600 1267.200 ;
        RECT 1.905 1263.120 798.495 1265.800 ;
        RECT 4.400 1261.720 795.600 1263.120 ;
        RECT 1.905 1259.040 798.495 1261.720 ;
        RECT 4.400 1257.640 795.600 1259.040 ;
        RECT 1.905 1254.960 798.495 1257.640 ;
        RECT 4.400 1253.560 795.600 1254.960 ;
        RECT 1.905 1250.880 798.495 1253.560 ;
        RECT 4.400 1249.480 795.600 1250.880 ;
        RECT 1.905 1246.800 798.495 1249.480 ;
        RECT 4.400 1245.400 795.600 1246.800 ;
        RECT 1.905 1242.720 798.495 1245.400 ;
        RECT 4.400 1241.320 795.600 1242.720 ;
        RECT 1.905 1238.640 798.495 1241.320 ;
        RECT 4.400 1237.240 795.600 1238.640 ;
        RECT 1.905 1234.560 798.495 1237.240 ;
        RECT 4.400 1233.160 795.600 1234.560 ;
        RECT 1.905 1230.480 798.495 1233.160 ;
        RECT 4.400 1229.080 795.600 1230.480 ;
        RECT 1.905 1226.400 798.495 1229.080 ;
        RECT 4.400 1225.000 795.600 1226.400 ;
        RECT 1.905 1222.320 798.495 1225.000 ;
        RECT 4.400 1220.920 795.600 1222.320 ;
        RECT 1.905 1218.240 798.495 1220.920 ;
        RECT 4.400 1216.840 795.600 1218.240 ;
        RECT 1.905 1214.160 798.495 1216.840 ;
        RECT 4.400 1212.760 795.600 1214.160 ;
        RECT 1.905 1210.080 798.495 1212.760 ;
        RECT 4.400 1208.680 795.600 1210.080 ;
        RECT 1.905 1206.000 798.495 1208.680 ;
        RECT 4.400 1204.600 795.600 1206.000 ;
        RECT 1.905 1201.920 798.495 1204.600 ;
        RECT 4.400 1200.520 795.600 1201.920 ;
        RECT 1.905 1197.840 798.495 1200.520 ;
        RECT 4.400 1196.440 795.600 1197.840 ;
        RECT 1.905 1193.760 798.495 1196.440 ;
        RECT 4.400 1192.360 795.600 1193.760 ;
        RECT 1.905 1189.680 798.495 1192.360 ;
        RECT 4.400 1188.280 795.600 1189.680 ;
        RECT 1.905 1185.600 798.495 1188.280 ;
        RECT 4.400 1184.200 795.600 1185.600 ;
        RECT 1.905 1181.520 798.495 1184.200 ;
        RECT 4.400 1180.120 795.600 1181.520 ;
        RECT 1.905 1177.440 798.495 1180.120 ;
        RECT 4.400 1176.040 795.600 1177.440 ;
        RECT 1.905 1173.360 798.495 1176.040 ;
        RECT 4.400 1171.960 795.600 1173.360 ;
        RECT 1.905 1169.280 798.495 1171.960 ;
        RECT 4.400 1167.880 795.600 1169.280 ;
        RECT 1.905 1165.200 798.495 1167.880 ;
        RECT 4.400 1163.800 795.600 1165.200 ;
        RECT 1.905 1161.120 798.495 1163.800 ;
        RECT 4.400 1159.720 795.600 1161.120 ;
        RECT 1.905 1157.040 798.495 1159.720 ;
        RECT 4.400 1155.640 795.600 1157.040 ;
        RECT 1.905 1152.960 798.495 1155.640 ;
        RECT 4.400 1151.560 795.600 1152.960 ;
        RECT 1.905 1148.880 798.495 1151.560 ;
        RECT 4.400 1147.480 795.600 1148.880 ;
        RECT 1.905 1144.800 798.495 1147.480 ;
        RECT 4.400 1143.400 795.600 1144.800 ;
        RECT 1.905 1140.720 798.495 1143.400 ;
        RECT 4.400 1139.320 795.600 1140.720 ;
        RECT 1.905 1136.640 798.495 1139.320 ;
        RECT 4.400 1135.240 795.600 1136.640 ;
        RECT 1.905 1132.560 798.495 1135.240 ;
        RECT 4.400 1131.160 795.600 1132.560 ;
        RECT 1.905 1128.480 798.495 1131.160 ;
        RECT 4.400 1127.080 795.600 1128.480 ;
        RECT 1.905 1124.400 798.495 1127.080 ;
        RECT 4.400 1123.000 795.600 1124.400 ;
        RECT 1.905 1120.320 798.495 1123.000 ;
        RECT 4.400 1118.920 795.600 1120.320 ;
        RECT 1.905 1116.240 798.495 1118.920 ;
        RECT 4.400 1114.840 795.600 1116.240 ;
        RECT 1.905 1112.160 798.495 1114.840 ;
        RECT 4.400 1110.760 795.600 1112.160 ;
        RECT 1.905 1108.080 798.495 1110.760 ;
        RECT 4.400 1106.680 795.600 1108.080 ;
        RECT 1.905 1104.000 798.495 1106.680 ;
        RECT 4.400 1102.600 795.600 1104.000 ;
        RECT 1.905 1099.920 798.495 1102.600 ;
        RECT 4.400 1098.520 795.600 1099.920 ;
        RECT 1.905 1095.840 798.495 1098.520 ;
        RECT 4.400 1094.440 795.600 1095.840 ;
        RECT 1.905 1091.760 798.495 1094.440 ;
        RECT 4.400 1090.360 795.600 1091.760 ;
        RECT 1.905 1087.680 798.495 1090.360 ;
        RECT 4.400 1086.280 795.600 1087.680 ;
        RECT 1.905 1083.600 798.495 1086.280 ;
        RECT 4.400 1082.200 795.600 1083.600 ;
        RECT 1.905 1079.520 798.495 1082.200 ;
        RECT 4.400 1078.120 795.600 1079.520 ;
        RECT 1.905 1075.440 798.495 1078.120 ;
        RECT 4.400 1074.040 795.600 1075.440 ;
        RECT 1.905 1071.360 798.495 1074.040 ;
        RECT 4.400 1069.960 795.600 1071.360 ;
        RECT 1.905 1067.280 798.495 1069.960 ;
        RECT 4.400 1065.880 795.600 1067.280 ;
        RECT 1.905 1063.200 798.495 1065.880 ;
        RECT 4.400 1061.800 795.600 1063.200 ;
        RECT 1.905 1059.120 798.495 1061.800 ;
        RECT 4.400 1057.720 795.600 1059.120 ;
        RECT 1.905 1055.040 798.495 1057.720 ;
        RECT 4.400 1053.640 795.600 1055.040 ;
        RECT 1.905 1050.960 798.495 1053.640 ;
        RECT 4.400 1049.560 795.600 1050.960 ;
        RECT 1.905 1046.880 798.495 1049.560 ;
        RECT 4.400 1045.480 795.600 1046.880 ;
        RECT 1.905 1042.800 798.495 1045.480 ;
        RECT 4.400 1041.400 795.600 1042.800 ;
        RECT 1.905 1038.720 798.495 1041.400 ;
        RECT 4.400 1037.320 795.600 1038.720 ;
        RECT 1.905 1034.640 798.495 1037.320 ;
        RECT 4.400 1033.240 795.600 1034.640 ;
        RECT 1.905 1030.560 798.495 1033.240 ;
        RECT 4.400 1029.160 795.600 1030.560 ;
        RECT 1.905 1026.480 798.495 1029.160 ;
        RECT 4.400 1025.080 795.600 1026.480 ;
        RECT 1.905 1022.400 798.495 1025.080 ;
        RECT 4.400 1021.000 795.600 1022.400 ;
        RECT 1.905 1018.320 798.495 1021.000 ;
        RECT 4.400 1016.920 795.600 1018.320 ;
        RECT 1.905 1014.240 798.495 1016.920 ;
        RECT 4.400 1012.840 795.600 1014.240 ;
        RECT 1.905 1010.160 798.495 1012.840 ;
        RECT 4.400 1008.760 795.600 1010.160 ;
        RECT 1.905 1006.080 798.495 1008.760 ;
        RECT 4.400 1004.680 795.600 1006.080 ;
        RECT 1.905 1002.000 798.495 1004.680 ;
        RECT 4.400 1000.600 795.600 1002.000 ;
        RECT 1.905 997.920 798.495 1000.600 ;
        RECT 4.400 996.520 795.600 997.920 ;
        RECT 1.905 993.840 798.495 996.520 ;
        RECT 4.400 992.440 795.600 993.840 ;
        RECT 1.905 989.760 798.495 992.440 ;
        RECT 4.400 988.360 795.600 989.760 ;
        RECT 1.905 985.680 798.495 988.360 ;
        RECT 4.400 984.280 795.600 985.680 ;
        RECT 1.905 981.600 798.495 984.280 ;
        RECT 4.400 980.200 795.600 981.600 ;
        RECT 1.905 977.520 798.495 980.200 ;
        RECT 4.400 976.120 795.600 977.520 ;
        RECT 1.905 973.440 798.495 976.120 ;
        RECT 4.400 972.040 795.600 973.440 ;
        RECT 1.905 969.360 798.495 972.040 ;
        RECT 4.400 967.960 795.600 969.360 ;
        RECT 1.905 965.280 798.495 967.960 ;
        RECT 4.400 963.880 795.600 965.280 ;
        RECT 1.905 961.200 798.495 963.880 ;
        RECT 4.400 959.800 795.600 961.200 ;
        RECT 1.905 957.120 798.495 959.800 ;
        RECT 4.400 955.720 795.600 957.120 ;
        RECT 1.905 953.040 798.495 955.720 ;
        RECT 4.400 951.640 795.600 953.040 ;
        RECT 1.905 948.960 798.495 951.640 ;
        RECT 4.400 947.560 795.600 948.960 ;
        RECT 1.905 944.880 798.495 947.560 ;
        RECT 4.400 943.480 795.600 944.880 ;
        RECT 1.905 940.800 798.495 943.480 ;
        RECT 4.400 939.400 795.600 940.800 ;
        RECT 1.905 936.720 798.495 939.400 ;
        RECT 4.400 935.320 795.600 936.720 ;
        RECT 1.905 932.640 798.495 935.320 ;
        RECT 4.400 931.240 795.600 932.640 ;
        RECT 1.905 928.560 798.495 931.240 ;
        RECT 4.400 927.160 795.600 928.560 ;
        RECT 1.905 924.480 798.495 927.160 ;
        RECT 4.400 923.080 795.600 924.480 ;
        RECT 1.905 920.400 798.495 923.080 ;
        RECT 4.400 919.000 795.600 920.400 ;
        RECT 1.905 916.320 798.495 919.000 ;
        RECT 4.400 914.920 795.600 916.320 ;
        RECT 1.905 912.240 798.495 914.920 ;
        RECT 4.400 910.840 795.600 912.240 ;
        RECT 1.905 908.160 798.495 910.840 ;
        RECT 4.400 906.760 795.600 908.160 ;
        RECT 1.905 904.080 798.495 906.760 ;
        RECT 4.400 902.680 795.600 904.080 ;
        RECT 1.905 900.000 798.495 902.680 ;
        RECT 4.400 898.600 795.600 900.000 ;
        RECT 1.905 895.920 798.495 898.600 ;
        RECT 4.400 894.520 795.600 895.920 ;
        RECT 1.905 891.840 798.495 894.520 ;
        RECT 4.400 890.440 795.600 891.840 ;
        RECT 1.905 887.760 798.495 890.440 ;
        RECT 4.400 886.360 795.600 887.760 ;
        RECT 1.905 883.680 798.495 886.360 ;
        RECT 4.400 882.280 795.600 883.680 ;
        RECT 1.905 879.600 798.495 882.280 ;
        RECT 4.400 878.200 795.600 879.600 ;
        RECT 1.905 875.520 798.495 878.200 ;
        RECT 4.400 874.120 795.600 875.520 ;
        RECT 1.905 871.440 798.495 874.120 ;
        RECT 4.400 870.040 795.600 871.440 ;
        RECT 1.905 867.360 798.495 870.040 ;
        RECT 4.400 865.960 795.600 867.360 ;
        RECT 1.905 863.280 798.495 865.960 ;
        RECT 4.400 861.880 795.600 863.280 ;
        RECT 1.905 859.200 798.495 861.880 ;
        RECT 4.400 857.800 795.600 859.200 ;
        RECT 1.905 855.120 798.495 857.800 ;
        RECT 4.400 853.720 795.600 855.120 ;
        RECT 1.905 851.040 798.495 853.720 ;
        RECT 4.400 849.640 795.600 851.040 ;
        RECT 1.905 846.960 798.495 849.640 ;
        RECT 4.400 845.560 795.600 846.960 ;
        RECT 1.905 842.880 798.495 845.560 ;
        RECT 4.400 841.480 795.600 842.880 ;
        RECT 1.905 838.800 798.495 841.480 ;
        RECT 4.400 837.400 795.600 838.800 ;
        RECT 1.905 834.720 798.495 837.400 ;
        RECT 4.400 833.320 795.600 834.720 ;
        RECT 1.905 830.640 798.495 833.320 ;
        RECT 4.400 829.240 795.600 830.640 ;
        RECT 1.905 826.560 798.495 829.240 ;
        RECT 4.400 825.160 795.600 826.560 ;
        RECT 1.905 822.480 798.495 825.160 ;
        RECT 4.400 821.080 795.600 822.480 ;
        RECT 1.905 818.400 798.495 821.080 ;
        RECT 4.400 817.000 795.600 818.400 ;
        RECT 1.905 814.320 798.495 817.000 ;
        RECT 4.400 812.920 795.600 814.320 ;
        RECT 1.905 810.240 798.495 812.920 ;
        RECT 4.400 808.840 795.600 810.240 ;
        RECT 1.905 806.160 798.495 808.840 ;
        RECT 4.400 804.760 795.600 806.160 ;
        RECT 1.905 802.080 798.495 804.760 ;
        RECT 4.400 800.680 795.600 802.080 ;
        RECT 1.905 798.000 798.495 800.680 ;
        RECT 4.400 796.600 795.600 798.000 ;
        RECT 1.905 793.920 798.495 796.600 ;
        RECT 4.400 792.520 795.600 793.920 ;
        RECT 1.905 789.840 798.495 792.520 ;
        RECT 4.400 788.440 795.600 789.840 ;
        RECT 1.905 785.760 798.495 788.440 ;
        RECT 4.400 784.360 795.600 785.760 ;
        RECT 1.905 781.680 798.495 784.360 ;
        RECT 4.400 780.280 795.600 781.680 ;
        RECT 1.905 777.600 798.495 780.280 ;
        RECT 4.400 776.200 795.600 777.600 ;
        RECT 1.905 773.520 798.495 776.200 ;
        RECT 4.400 772.120 795.600 773.520 ;
        RECT 1.905 769.440 798.495 772.120 ;
        RECT 4.400 768.040 795.600 769.440 ;
        RECT 1.905 765.360 798.495 768.040 ;
        RECT 4.400 763.960 795.600 765.360 ;
        RECT 1.905 761.280 798.495 763.960 ;
        RECT 4.400 759.880 795.600 761.280 ;
        RECT 1.905 757.200 798.495 759.880 ;
        RECT 4.400 755.800 795.600 757.200 ;
        RECT 1.905 753.120 798.495 755.800 ;
        RECT 4.400 751.720 795.600 753.120 ;
        RECT 1.905 749.040 798.495 751.720 ;
        RECT 4.400 747.640 795.600 749.040 ;
        RECT 1.905 744.960 798.495 747.640 ;
        RECT 4.400 743.560 795.600 744.960 ;
        RECT 1.905 740.880 798.495 743.560 ;
        RECT 4.400 739.480 795.600 740.880 ;
        RECT 1.905 736.800 798.495 739.480 ;
        RECT 4.400 735.400 795.600 736.800 ;
        RECT 1.905 732.720 798.495 735.400 ;
        RECT 4.400 731.320 795.600 732.720 ;
        RECT 1.905 728.640 798.495 731.320 ;
        RECT 4.400 727.240 795.600 728.640 ;
        RECT 1.905 724.560 798.495 727.240 ;
        RECT 4.400 723.160 795.600 724.560 ;
        RECT 1.905 720.480 798.495 723.160 ;
        RECT 4.400 719.080 795.600 720.480 ;
        RECT 1.905 716.400 798.495 719.080 ;
        RECT 4.400 715.000 795.600 716.400 ;
        RECT 1.905 712.320 798.495 715.000 ;
        RECT 4.400 710.920 795.600 712.320 ;
        RECT 1.905 708.240 798.495 710.920 ;
        RECT 4.400 706.840 795.600 708.240 ;
        RECT 1.905 704.160 798.495 706.840 ;
        RECT 4.400 702.760 795.600 704.160 ;
        RECT 1.905 700.080 798.495 702.760 ;
        RECT 4.400 698.680 795.600 700.080 ;
        RECT 1.905 696.000 798.495 698.680 ;
        RECT 4.400 694.600 795.600 696.000 ;
        RECT 1.905 691.920 798.495 694.600 ;
        RECT 4.400 690.520 795.600 691.920 ;
        RECT 1.905 687.840 798.495 690.520 ;
        RECT 4.400 686.440 795.600 687.840 ;
        RECT 1.905 683.760 798.495 686.440 ;
        RECT 4.400 682.360 795.600 683.760 ;
        RECT 1.905 679.680 798.495 682.360 ;
        RECT 4.400 678.280 795.600 679.680 ;
        RECT 1.905 675.600 798.495 678.280 ;
        RECT 4.400 674.200 795.600 675.600 ;
        RECT 1.905 671.520 798.495 674.200 ;
        RECT 4.400 670.120 795.600 671.520 ;
        RECT 1.905 667.440 798.495 670.120 ;
        RECT 4.400 666.040 795.600 667.440 ;
        RECT 1.905 663.360 798.495 666.040 ;
        RECT 4.400 661.960 795.600 663.360 ;
        RECT 1.905 659.280 798.495 661.960 ;
        RECT 4.400 657.880 795.600 659.280 ;
        RECT 1.905 655.200 798.495 657.880 ;
        RECT 4.400 653.800 795.600 655.200 ;
        RECT 1.905 651.120 798.495 653.800 ;
        RECT 4.400 649.720 795.600 651.120 ;
        RECT 1.905 647.040 798.495 649.720 ;
        RECT 4.400 645.640 795.600 647.040 ;
        RECT 1.905 642.960 798.495 645.640 ;
        RECT 4.400 641.560 795.600 642.960 ;
        RECT 1.905 638.880 798.495 641.560 ;
        RECT 4.400 637.480 795.600 638.880 ;
        RECT 1.905 634.800 798.495 637.480 ;
        RECT 4.400 633.400 795.600 634.800 ;
        RECT 1.905 630.720 798.495 633.400 ;
        RECT 4.400 629.320 795.600 630.720 ;
        RECT 1.905 626.640 798.495 629.320 ;
        RECT 4.400 625.240 795.600 626.640 ;
        RECT 1.905 622.560 798.495 625.240 ;
        RECT 4.400 621.160 795.600 622.560 ;
        RECT 1.905 618.480 798.495 621.160 ;
        RECT 4.400 617.080 795.600 618.480 ;
        RECT 1.905 614.400 798.495 617.080 ;
        RECT 4.400 613.000 795.600 614.400 ;
        RECT 1.905 610.320 798.495 613.000 ;
        RECT 4.400 608.920 795.600 610.320 ;
        RECT 1.905 606.240 798.495 608.920 ;
        RECT 4.400 604.840 795.600 606.240 ;
        RECT 1.905 602.160 798.495 604.840 ;
        RECT 4.400 600.760 795.600 602.160 ;
        RECT 1.905 598.080 798.495 600.760 ;
        RECT 4.400 596.680 795.600 598.080 ;
        RECT 1.905 594.000 798.495 596.680 ;
        RECT 4.400 592.600 795.600 594.000 ;
        RECT 1.905 589.920 798.495 592.600 ;
        RECT 4.400 588.520 795.600 589.920 ;
        RECT 1.905 585.840 798.495 588.520 ;
        RECT 4.400 584.440 795.600 585.840 ;
        RECT 1.905 581.760 798.495 584.440 ;
        RECT 4.400 580.360 795.600 581.760 ;
        RECT 1.905 577.680 798.495 580.360 ;
        RECT 4.400 576.280 795.600 577.680 ;
        RECT 1.905 573.600 798.495 576.280 ;
        RECT 4.400 572.200 795.600 573.600 ;
        RECT 1.905 569.520 798.495 572.200 ;
        RECT 4.400 568.120 795.600 569.520 ;
        RECT 1.905 565.440 798.495 568.120 ;
        RECT 4.400 564.040 795.600 565.440 ;
        RECT 1.905 561.360 798.495 564.040 ;
        RECT 4.400 559.960 795.600 561.360 ;
        RECT 1.905 557.280 798.495 559.960 ;
        RECT 4.400 555.880 795.600 557.280 ;
        RECT 1.905 553.200 798.495 555.880 ;
        RECT 4.400 551.800 795.600 553.200 ;
        RECT 1.905 549.120 798.495 551.800 ;
        RECT 4.400 547.720 795.600 549.120 ;
        RECT 1.905 545.040 798.495 547.720 ;
        RECT 4.400 543.640 795.600 545.040 ;
        RECT 1.905 540.960 798.495 543.640 ;
        RECT 4.400 539.560 795.600 540.960 ;
        RECT 1.905 536.880 798.495 539.560 ;
        RECT 4.400 535.480 795.600 536.880 ;
        RECT 1.905 532.800 798.495 535.480 ;
        RECT 4.400 531.400 795.600 532.800 ;
        RECT 1.905 528.720 798.495 531.400 ;
        RECT 4.400 527.320 795.600 528.720 ;
        RECT 1.905 524.640 798.495 527.320 ;
        RECT 4.400 523.240 795.600 524.640 ;
        RECT 1.905 520.560 798.495 523.240 ;
        RECT 4.400 519.160 795.600 520.560 ;
        RECT 1.905 516.480 798.495 519.160 ;
        RECT 4.400 515.080 795.600 516.480 ;
        RECT 1.905 512.400 798.495 515.080 ;
        RECT 4.400 511.000 795.600 512.400 ;
        RECT 1.905 508.320 798.495 511.000 ;
        RECT 4.400 506.920 795.600 508.320 ;
        RECT 1.905 504.240 798.495 506.920 ;
        RECT 4.400 502.840 795.600 504.240 ;
        RECT 1.905 500.160 798.495 502.840 ;
        RECT 4.400 498.760 795.600 500.160 ;
        RECT 1.905 496.080 798.495 498.760 ;
        RECT 4.400 494.680 795.600 496.080 ;
        RECT 1.905 492.000 798.495 494.680 ;
        RECT 4.400 490.600 795.600 492.000 ;
        RECT 1.905 487.920 798.495 490.600 ;
        RECT 4.400 486.520 795.600 487.920 ;
        RECT 1.905 483.840 798.495 486.520 ;
        RECT 4.400 482.440 795.600 483.840 ;
        RECT 1.905 479.760 798.495 482.440 ;
        RECT 4.400 478.360 795.600 479.760 ;
        RECT 1.905 475.680 798.495 478.360 ;
        RECT 4.400 474.280 795.600 475.680 ;
        RECT 1.905 471.600 798.495 474.280 ;
        RECT 4.400 470.200 795.600 471.600 ;
        RECT 1.905 467.520 798.495 470.200 ;
        RECT 4.400 466.120 795.600 467.520 ;
        RECT 1.905 463.440 798.495 466.120 ;
        RECT 4.400 462.040 795.600 463.440 ;
        RECT 1.905 459.360 798.495 462.040 ;
        RECT 4.400 457.960 795.600 459.360 ;
        RECT 1.905 455.280 798.495 457.960 ;
        RECT 4.400 453.880 795.600 455.280 ;
        RECT 1.905 451.200 798.495 453.880 ;
        RECT 4.400 449.800 795.600 451.200 ;
        RECT 1.905 447.120 798.495 449.800 ;
        RECT 4.400 445.720 795.600 447.120 ;
        RECT 1.905 443.040 798.495 445.720 ;
        RECT 4.400 441.640 795.600 443.040 ;
        RECT 1.905 438.960 798.495 441.640 ;
        RECT 4.400 437.560 795.600 438.960 ;
        RECT 1.905 434.880 798.495 437.560 ;
        RECT 4.400 433.480 795.600 434.880 ;
        RECT 1.905 430.800 798.495 433.480 ;
        RECT 4.400 429.400 795.600 430.800 ;
        RECT 1.905 426.720 798.495 429.400 ;
        RECT 4.400 425.320 795.600 426.720 ;
        RECT 1.905 422.640 798.495 425.320 ;
        RECT 4.400 421.240 795.600 422.640 ;
        RECT 1.905 418.560 798.495 421.240 ;
        RECT 4.400 417.160 795.600 418.560 ;
        RECT 1.905 414.480 798.495 417.160 ;
        RECT 4.400 413.080 795.600 414.480 ;
        RECT 1.905 410.400 798.495 413.080 ;
        RECT 4.400 409.000 795.600 410.400 ;
        RECT 1.905 406.320 798.495 409.000 ;
        RECT 4.400 404.920 795.600 406.320 ;
        RECT 1.905 402.240 798.495 404.920 ;
        RECT 4.400 400.840 795.600 402.240 ;
        RECT 1.905 398.160 798.495 400.840 ;
        RECT 4.400 396.760 795.600 398.160 ;
        RECT 1.905 394.080 798.495 396.760 ;
        RECT 4.400 392.680 795.600 394.080 ;
        RECT 1.905 390.000 798.495 392.680 ;
        RECT 4.400 388.600 795.600 390.000 ;
        RECT 1.905 385.920 798.495 388.600 ;
        RECT 4.400 384.520 795.600 385.920 ;
        RECT 1.905 381.840 798.495 384.520 ;
        RECT 4.400 380.440 795.600 381.840 ;
        RECT 1.905 377.760 798.495 380.440 ;
        RECT 4.400 376.360 795.600 377.760 ;
        RECT 1.905 373.680 798.495 376.360 ;
        RECT 4.400 372.280 795.600 373.680 ;
        RECT 1.905 369.600 798.495 372.280 ;
        RECT 4.400 368.200 795.600 369.600 ;
        RECT 1.905 365.520 798.495 368.200 ;
        RECT 4.400 364.120 795.600 365.520 ;
        RECT 1.905 361.440 798.495 364.120 ;
        RECT 4.400 360.040 795.600 361.440 ;
        RECT 1.905 357.360 798.495 360.040 ;
        RECT 4.400 355.960 795.600 357.360 ;
        RECT 1.905 353.280 798.495 355.960 ;
        RECT 4.400 351.880 795.600 353.280 ;
        RECT 1.905 349.200 798.495 351.880 ;
        RECT 4.400 347.800 795.600 349.200 ;
        RECT 1.905 345.120 798.495 347.800 ;
        RECT 4.400 343.720 795.600 345.120 ;
        RECT 1.905 341.040 798.495 343.720 ;
        RECT 4.400 339.640 795.600 341.040 ;
        RECT 1.905 336.960 798.495 339.640 ;
        RECT 4.400 335.560 795.600 336.960 ;
        RECT 1.905 332.880 798.495 335.560 ;
        RECT 4.400 331.480 795.600 332.880 ;
        RECT 1.905 328.800 798.495 331.480 ;
        RECT 4.400 327.400 795.600 328.800 ;
        RECT 1.905 324.720 798.495 327.400 ;
        RECT 4.400 323.320 795.600 324.720 ;
        RECT 1.905 320.640 798.495 323.320 ;
        RECT 4.400 319.240 795.600 320.640 ;
        RECT 1.905 316.560 798.495 319.240 ;
        RECT 4.400 315.160 795.600 316.560 ;
        RECT 1.905 312.480 798.495 315.160 ;
        RECT 4.400 311.080 795.600 312.480 ;
        RECT 1.905 308.400 798.495 311.080 ;
        RECT 4.400 307.000 795.600 308.400 ;
        RECT 1.905 304.320 798.495 307.000 ;
        RECT 4.400 302.920 795.600 304.320 ;
        RECT 1.905 300.240 798.495 302.920 ;
        RECT 4.400 298.840 795.600 300.240 ;
        RECT 1.905 296.160 798.495 298.840 ;
        RECT 4.400 294.760 795.600 296.160 ;
        RECT 1.905 292.080 798.495 294.760 ;
        RECT 4.400 290.680 795.600 292.080 ;
        RECT 1.905 288.000 798.495 290.680 ;
        RECT 4.400 286.600 795.600 288.000 ;
        RECT 1.905 283.920 798.495 286.600 ;
        RECT 4.400 282.520 795.600 283.920 ;
        RECT 1.905 279.840 798.495 282.520 ;
        RECT 4.400 278.440 795.600 279.840 ;
        RECT 1.905 275.760 798.495 278.440 ;
        RECT 4.400 274.360 795.600 275.760 ;
        RECT 1.905 271.680 798.495 274.360 ;
        RECT 4.400 270.280 795.600 271.680 ;
        RECT 1.905 267.600 798.495 270.280 ;
        RECT 4.400 266.200 795.600 267.600 ;
        RECT 1.905 263.520 798.495 266.200 ;
        RECT 4.400 262.120 795.600 263.520 ;
        RECT 1.905 259.440 798.495 262.120 ;
        RECT 4.400 258.040 795.600 259.440 ;
        RECT 1.905 255.360 798.495 258.040 ;
        RECT 4.400 253.960 795.600 255.360 ;
        RECT 1.905 251.280 798.495 253.960 ;
        RECT 4.400 249.880 795.600 251.280 ;
        RECT 1.905 247.200 798.495 249.880 ;
        RECT 4.400 245.800 795.600 247.200 ;
        RECT 1.905 243.120 798.495 245.800 ;
        RECT 4.400 241.720 795.600 243.120 ;
        RECT 1.905 239.040 798.495 241.720 ;
        RECT 4.400 237.640 795.600 239.040 ;
        RECT 1.905 234.960 798.495 237.640 ;
        RECT 4.400 233.560 795.600 234.960 ;
        RECT 1.905 230.880 798.495 233.560 ;
        RECT 4.400 229.480 795.600 230.880 ;
        RECT 1.905 226.800 798.495 229.480 ;
        RECT 4.400 225.400 795.600 226.800 ;
        RECT 1.905 222.720 798.495 225.400 ;
        RECT 4.400 221.320 795.600 222.720 ;
        RECT 1.905 218.640 798.495 221.320 ;
        RECT 4.400 217.240 795.600 218.640 ;
        RECT 1.905 214.560 798.495 217.240 ;
        RECT 4.400 213.160 795.600 214.560 ;
        RECT 1.905 210.480 798.495 213.160 ;
        RECT 4.400 209.080 795.600 210.480 ;
        RECT 1.905 206.400 798.495 209.080 ;
        RECT 4.400 205.000 795.600 206.400 ;
        RECT 1.905 202.320 798.495 205.000 ;
        RECT 4.400 200.920 795.600 202.320 ;
        RECT 1.905 198.240 798.495 200.920 ;
        RECT 4.400 196.840 795.600 198.240 ;
        RECT 1.905 194.160 798.495 196.840 ;
        RECT 4.400 192.760 795.600 194.160 ;
        RECT 1.905 190.080 798.495 192.760 ;
        RECT 4.400 188.680 795.600 190.080 ;
        RECT 1.905 186.000 798.495 188.680 ;
        RECT 4.400 184.600 795.600 186.000 ;
        RECT 1.905 181.920 798.495 184.600 ;
        RECT 4.400 180.520 795.600 181.920 ;
        RECT 1.905 177.840 798.495 180.520 ;
        RECT 4.400 176.440 795.600 177.840 ;
        RECT 1.905 173.760 798.495 176.440 ;
        RECT 4.400 172.360 795.600 173.760 ;
        RECT 1.905 169.680 798.495 172.360 ;
        RECT 4.400 168.280 795.600 169.680 ;
        RECT 1.905 165.600 798.495 168.280 ;
        RECT 4.400 164.200 795.600 165.600 ;
        RECT 1.905 161.520 798.495 164.200 ;
        RECT 4.400 160.120 795.600 161.520 ;
        RECT 1.905 157.440 798.495 160.120 ;
        RECT 4.400 156.040 795.600 157.440 ;
        RECT 1.905 10.715 798.495 156.040 ;
      LAYER met4 ;
        RECT 3.055 162.015 20.640 2386.625 ;
        RECT 23.040 162.015 97.440 2386.625 ;
        RECT 99.840 162.015 174.240 2386.625 ;
        RECT 176.640 162.015 251.040 2386.625 ;
        RECT 253.440 162.015 327.840 2386.625 ;
        RECT 330.240 162.015 404.640 2386.625 ;
        RECT 407.040 162.015 481.440 2386.625 ;
        RECT 483.840 162.015 558.240 2386.625 ;
        RECT 560.640 162.015 635.040 2386.625 ;
        RECT 637.440 162.015 711.840 2386.625 ;
        RECT 714.240 162.015 783.545 2386.625 ;
  END
END IMPACTSram
END LIBRARY

