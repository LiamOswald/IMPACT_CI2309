VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO IMPACTSram
  CLASS BLOCK ;
  FOREIGN IMPACTSram ;
  ORIGIN 0.790 43.350 ;
  SIZE 221.940 BY 62.720 ;
  PIN BL0
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER li1 ;
        RECT 1.420 14.860 1.870 15.310 ;
        RECT 1.420 11.250 1.870 11.700 ;
        RECT 1.420 7.640 1.870 8.090 ;
        RECT 1.420 4.030 1.870 4.480 ;
        RECT 1.420 0.420 1.870 0.870 ;
        RECT 1.420 -3.190 1.870 -2.740 ;
        RECT 1.420 -6.800 1.870 -6.350 ;
        RECT 1.420 -10.410 1.870 -9.960 ;
        RECT 1.420 -14.020 1.870 -13.570 ;
        RECT 1.420 -17.630 1.870 -17.180 ;
        RECT 1.420 -21.240 1.870 -20.790 ;
        RECT 1.420 -24.850 1.870 -24.400 ;
        RECT 1.420 -28.460 1.870 -28.010 ;
        RECT 1.420 -32.070 1.870 -31.620 ;
        RECT 1.420 -35.680 1.870 -35.230 ;
        RECT 1.420 -39.290 1.870 -38.840 ;
      LAYER mcon ;
        RECT 1.520 14.960 1.770 15.210 ;
        RECT 1.520 11.350 1.770 11.600 ;
        RECT 1.520 7.740 1.770 7.990 ;
        RECT 1.520 4.130 1.770 4.380 ;
        RECT 1.520 0.520 1.770 0.770 ;
        RECT 1.520 -3.090 1.770 -2.840 ;
        RECT 1.520 -6.700 1.770 -6.450 ;
        RECT 1.520 -10.310 1.770 -10.060 ;
        RECT 1.520 -13.920 1.770 -13.670 ;
        RECT 1.520 -17.530 1.770 -17.280 ;
        RECT 1.520 -21.140 1.770 -20.890 ;
        RECT 1.520 -24.750 1.770 -24.500 ;
        RECT 1.520 -28.360 1.770 -28.110 ;
        RECT 1.520 -31.970 1.770 -31.720 ;
        RECT 1.520 -35.580 1.770 -35.330 ;
        RECT 1.520 -39.190 1.770 -38.940 ;
      LAYER met1 ;
        RECT 1.300 -43.100 1.980 19.120 ;
    END
  END BL0
  PIN BLb0
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER li1 ;
        RECT 6.520 16.660 6.970 17.110 ;
        RECT 6.520 13.050 6.970 13.510 ;
        RECT 6.520 9.440 6.970 9.900 ;
        RECT 6.520 5.830 6.970 6.290 ;
        RECT 6.520 2.220 6.970 2.680 ;
        RECT 6.520 -1.390 6.970 -0.930 ;
        RECT 6.520 -5.000 6.970 -4.540 ;
        RECT 6.520 -8.610 6.970 -8.150 ;
        RECT 6.520 -12.220 6.970 -11.760 ;
        RECT 6.520 -15.830 6.970 -15.370 ;
        RECT 6.520 -19.440 6.970 -18.980 ;
        RECT 6.520 -23.050 6.970 -22.590 ;
        RECT 6.520 -26.660 6.970 -26.200 ;
        RECT 6.520 -30.270 6.970 -29.810 ;
        RECT 6.520 -33.880 6.970 -33.420 ;
        RECT 6.520 -37.490 6.970 -37.030 ;
        RECT 6.520 -41.090 6.970 -40.640 ;
      LAYER mcon ;
        RECT 6.620 16.760 6.880 17.020 ;
        RECT 6.620 13.150 6.880 13.410 ;
        RECT 6.620 9.540 6.880 9.800 ;
        RECT 6.620 5.930 6.880 6.190 ;
        RECT 6.620 2.320 6.880 2.580 ;
        RECT 6.620 -1.290 6.880 -1.030 ;
        RECT 6.620 -4.900 6.880 -4.640 ;
        RECT 6.620 -8.510 6.880 -8.250 ;
        RECT 6.620 -12.120 6.880 -11.860 ;
        RECT 6.620 -15.730 6.880 -15.470 ;
        RECT 6.620 -19.340 6.880 -19.080 ;
        RECT 6.620 -22.950 6.880 -22.690 ;
        RECT 6.620 -26.560 6.880 -26.300 ;
        RECT 6.620 -30.170 6.880 -29.910 ;
        RECT 6.620 -33.780 6.880 -33.520 ;
        RECT 6.620 -37.390 6.880 -37.130 ;
        RECT 6.620 -41.000 6.880 -40.740 ;
      LAYER met1 ;
        RECT 6.400 -43.120 7.080 19.140 ;
    END
  END BLb0
  PIN BL1
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER li1 ;
        RECT 8.160 16.660 8.610 17.110 ;
        RECT 8.160 13.050 8.610 13.510 ;
        RECT 8.160 9.440 8.610 9.900 ;
        RECT 8.160 5.830 8.610 6.290 ;
        RECT 8.160 2.220 8.610 2.680 ;
        RECT 8.160 -1.390 8.610 -0.930 ;
        RECT 8.160 -5.000 8.610 -4.540 ;
        RECT 8.160 -8.610 8.610 -8.150 ;
        RECT 8.160 -12.220 8.610 -11.760 ;
        RECT 8.160 -15.830 8.610 -15.370 ;
        RECT 8.160 -19.440 8.610 -18.980 ;
        RECT 8.160 -23.050 8.610 -22.590 ;
        RECT 8.160 -26.660 8.610 -26.200 ;
        RECT 8.160 -30.270 8.610 -29.810 ;
        RECT 8.160 -33.880 8.610 -33.420 ;
        RECT 8.160 -37.490 8.610 -37.030 ;
        RECT 8.160 -41.090 8.610 -40.640 ;
      LAYER mcon ;
        RECT 8.250 16.760 8.510 17.020 ;
        RECT 8.250 13.150 8.510 13.410 ;
        RECT 8.250 9.540 8.510 9.800 ;
        RECT 8.250 5.930 8.510 6.190 ;
        RECT 8.250 2.320 8.510 2.580 ;
        RECT 8.250 -1.290 8.510 -1.030 ;
        RECT 8.250 -4.900 8.510 -4.640 ;
        RECT 8.250 -8.510 8.510 -8.250 ;
        RECT 8.250 -12.120 8.510 -11.860 ;
        RECT 8.250 -15.730 8.510 -15.470 ;
        RECT 8.250 -19.340 8.510 -19.080 ;
        RECT 8.250 -22.950 8.510 -22.690 ;
        RECT 8.250 -26.560 8.510 -26.300 ;
        RECT 8.250 -30.170 8.510 -29.910 ;
        RECT 8.250 -33.780 8.510 -33.520 ;
        RECT 8.250 -37.390 8.510 -37.130 ;
        RECT 8.250 -41.000 8.510 -40.740 ;
      LAYER met1 ;
        RECT 8.040 -43.110 8.720 19.130 ;
    END
  END BL1
  PIN BLb1
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER li1 ;
        RECT 13.260 14.860 13.710 15.310 ;
        RECT 13.260 11.250 13.710 11.700 ;
        RECT 13.260 7.640 13.710 8.090 ;
        RECT 13.260 4.030 13.710 4.480 ;
        RECT 13.260 0.420 13.710 0.870 ;
        RECT 13.260 -3.190 13.710 -2.740 ;
        RECT 13.260 -6.800 13.710 -6.350 ;
        RECT 13.260 -10.410 13.710 -9.960 ;
        RECT 13.260 -14.020 13.710 -13.570 ;
        RECT 13.260 -17.630 13.710 -17.180 ;
        RECT 13.260 -21.240 13.710 -20.790 ;
        RECT 13.260 -24.850 13.710 -24.400 ;
        RECT 13.260 -28.460 13.710 -28.010 ;
        RECT 13.260 -32.070 13.710 -31.620 ;
        RECT 13.260 -35.680 13.710 -35.230 ;
        RECT 13.260 -39.290 13.710 -38.840 ;
      LAYER mcon ;
        RECT 13.360 14.960 13.610 15.210 ;
        RECT 13.360 11.350 13.610 11.600 ;
        RECT 13.360 7.740 13.610 7.990 ;
        RECT 13.360 4.130 13.610 4.380 ;
        RECT 13.360 0.520 13.610 0.770 ;
        RECT 13.360 -3.090 13.610 -2.840 ;
        RECT 13.360 -6.700 13.610 -6.450 ;
        RECT 13.360 -10.310 13.610 -10.060 ;
        RECT 13.360 -13.920 13.610 -13.670 ;
        RECT 13.360 -17.530 13.610 -17.280 ;
        RECT 13.360 -21.140 13.610 -20.890 ;
        RECT 13.360 -24.750 13.610 -24.500 ;
        RECT 13.360 -28.360 13.610 -28.110 ;
        RECT 13.360 -31.970 13.610 -31.720 ;
        RECT 13.360 -35.580 13.610 -35.330 ;
        RECT 13.360 -39.190 13.610 -38.940 ;
      LAYER met1 ;
        RECT 13.160 -43.110 13.840 19.130 ;
    END
  END BLb1
  PIN BL2
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER li1 ;
        RECT 14.920 14.860 15.370 15.310 ;
        RECT 14.920 11.250 15.370 11.700 ;
        RECT 14.920 7.640 15.370 8.090 ;
        RECT 14.920 4.030 15.370 4.480 ;
        RECT 14.920 0.420 15.370 0.870 ;
        RECT 14.920 -3.190 15.370 -2.740 ;
        RECT 14.920 -6.800 15.370 -6.350 ;
        RECT 14.920 -10.410 15.370 -9.960 ;
        RECT 14.920 -14.020 15.370 -13.570 ;
        RECT 14.920 -17.630 15.370 -17.180 ;
        RECT 14.920 -21.240 15.370 -20.790 ;
        RECT 14.920 -24.850 15.370 -24.400 ;
        RECT 14.920 -28.460 15.370 -28.010 ;
        RECT 14.920 -32.070 15.370 -31.620 ;
        RECT 14.920 -35.680 15.370 -35.230 ;
        RECT 14.920 -39.290 15.370 -38.840 ;
      LAYER mcon ;
        RECT 15.020 14.960 15.270 15.210 ;
        RECT 15.020 11.350 15.270 11.600 ;
        RECT 15.020 7.740 15.270 7.990 ;
        RECT 15.020 4.130 15.270 4.380 ;
        RECT 15.020 0.520 15.270 0.770 ;
        RECT 15.020 -3.090 15.270 -2.840 ;
        RECT 15.020 -6.700 15.270 -6.450 ;
        RECT 15.020 -10.310 15.270 -10.060 ;
        RECT 15.020 -13.920 15.270 -13.670 ;
        RECT 15.020 -17.530 15.270 -17.280 ;
        RECT 15.020 -21.140 15.270 -20.890 ;
        RECT 15.020 -24.750 15.270 -24.500 ;
        RECT 15.020 -28.360 15.270 -28.110 ;
        RECT 15.020 -31.970 15.270 -31.720 ;
        RECT 15.020 -35.580 15.270 -35.330 ;
        RECT 15.020 -39.190 15.270 -38.940 ;
      LAYER met1 ;
        RECT 14.800 -43.110 15.480 19.130 ;
    END
  END BL2
  PIN BLb2
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER li1 ;
        RECT 20.020 16.660 20.470 17.110 ;
        RECT 20.020 13.050 20.470 13.510 ;
        RECT 20.020 9.440 20.470 9.900 ;
        RECT 20.020 5.830 20.470 6.290 ;
        RECT 20.020 2.220 20.470 2.680 ;
        RECT 20.020 -1.390 20.470 -0.930 ;
        RECT 20.020 -5.000 20.470 -4.540 ;
        RECT 20.020 -8.610 20.470 -8.150 ;
        RECT 20.020 -12.220 20.470 -11.760 ;
        RECT 20.020 -15.830 20.470 -15.370 ;
        RECT 20.020 -19.440 20.470 -18.980 ;
        RECT 20.020 -23.050 20.470 -22.590 ;
        RECT 20.020 -26.660 20.470 -26.200 ;
        RECT 20.020 -30.270 20.470 -29.810 ;
        RECT 20.020 -33.880 20.470 -33.420 ;
        RECT 20.020 -37.490 20.470 -37.030 ;
        RECT 20.020 -41.090 20.470 -40.640 ;
      LAYER mcon ;
        RECT 20.120 16.760 20.380 17.020 ;
        RECT 20.120 13.150 20.380 13.410 ;
        RECT 20.120 9.540 20.380 9.800 ;
        RECT 20.120 5.930 20.380 6.190 ;
        RECT 20.120 2.320 20.380 2.580 ;
        RECT 20.120 -1.290 20.380 -1.030 ;
        RECT 20.120 -4.900 20.380 -4.640 ;
        RECT 20.120 -8.510 20.380 -8.250 ;
        RECT 20.120 -12.120 20.380 -11.860 ;
        RECT 20.120 -15.730 20.380 -15.470 ;
        RECT 20.120 -19.340 20.380 -19.080 ;
        RECT 20.120 -22.950 20.380 -22.690 ;
        RECT 20.120 -26.560 20.380 -26.300 ;
        RECT 20.120 -30.170 20.380 -29.910 ;
        RECT 20.120 -33.780 20.380 -33.520 ;
        RECT 20.120 -37.390 20.380 -37.130 ;
        RECT 20.120 -41.000 20.380 -40.740 ;
      LAYER met1 ;
        RECT 19.910 -43.120 20.590 19.140 ;
    END
  END BLb2
  PIN BL3
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER li1 ;
        RECT 21.660 16.660 22.110 17.110 ;
        RECT 21.660 13.050 22.110 13.510 ;
        RECT 21.660 9.440 22.110 9.900 ;
        RECT 21.660 5.830 22.110 6.290 ;
        RECT 21.660 2.220 22.110 2.680 ;
        RECT 21.660 -1.390 22.110 -0.930 ;
        RECT 21.660 -5.000 22.110 -4.540 ;
        RECT 21.660 -8.610 22.110 -8.150 ;
        RECT 21.660 -12.220 22.110 -11.760 ;
        RECT 21.660 -15.830 22.110 -15.370 ;
        RECT 21.660 -19.440 22.110 -18.980 ;
        RECT 21.660 -23.050 22.110 -22.590 ;
        RECT 21.660 -26.660 22.110 -26.200 ;
        RECT 21.660 -30.270 22.110 -29.810 ;
        RECT 21.660 -33.880 22.110 -33.420 ;
        RECT 21.660 -37.490 22.110 -37.030 ;
        RECT 21.660 -41.090 22.110 -40.640 ;
      LAYER mcon ;
        RECT 21.750 16.760 22.010 17.020 ;
        RECT 21.750 13.150 22.010 13.410 ;
        RECT 21.750 9.540 22.010 9.800 ;
        RECT 21.750 5.930 22.010 6.190 ;
        RECT 21.750 2.320 22.010 2.580 ;
        RECT 21.750 -1.290 22.010 -1.030 ;
        RECT 21.750 -4.900 22.010 -4.640 ;
        RECT 21.750 -8.510 22.010 -8.250 ;
        RECT 21.750 -12.120 22.010 -11.860 ;
        RECT 21.750 -15.730 22.010 -15.470 ;
        RECT 21.750 -19.340 22.010 -19.080 ;
        RECT 21.750 -22.950 22.010 -22.690 ;
        RECT 21.750 -26.560 22.010 -26.300 ;
        RECT 21.750 -30.170 22.010 -29.910 ;
        RECT 21.750 -33.780 22.010 -33.520 ;
        RECT 21.750 -37.390 22.010 -37.130 ;
        RECT 21.750 -41.000 22.010 -40.740 ;
      LAYER met1 ;
        RECT 21.550 -43.110 22.230 19.130 ;
    END
  END BL3
  PIN BLb3
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER li1 ;
        RECT 26.760 14.860 27.210 15.310 ;
        RECT 26.760 11.250 27.210 11.700 ;
        RECT 26.760 7.640 27.210 8.090 ;
        RECT 26.760 4.030 27.210 4.480 ;
        RECT 26.760 0.420 27.210 0.870 ;
        RECT 26.760 -3.190 27.210 -2.740 ;
        RECT 26.760 -6.800 27.210 -6.350 ;
        RECT 26.760 -10.410 27.210 -9.960 ;
        RECT 26.760 -14.020 27.210 -13.570 ;
        RECT 26.760 -17.630 27.210 -17.180 ;
        RECT 26.760 -21.240 27.210 -20.790 ;
        RECT 26.760 -24.850 27.210 -24.400 ;
        RECT 26.760 -28.460 27.210 -28.010 ;
        RECT 26.760 -32.070 27.210 -31.620 ;
        RECT 26.760 -35.680 27.210 -35.230 ;
        RECT 26.760 -39.290 27.210 -38.840 ;
      LAYER mcon ;
        RECT 26.860 14.960 27.110 15.210 ;
        RECT 26.860 11.350 27.110 11.600 ;
        RECT 26.860 7.740 27.110 7.990 ;
        RECT 26.860 4.130 27.110 4.380 ;
        RECT 26.860 0.520 27.110 0.770 ;
        RECT 26.860 -3.090 27.110 -2.840 ;
        RECT 26.860 -6.700 27.110 -6.450 ;
        RECT 26.860 -10.310 27.110 -10.060 ;
        RECT 26.860 -13.920 27.110 -13.670 ;
        RECT 26.860 -17.530 27.110 -17.280 ;
        RECT 26.860 -21.140 27.110 -20.890 ;
        RECT 26.860 -24.750 27.110 -24.500 ;
        RECT 26.860 -28.360 27.110 -28.110 ;
        RECT 26.860 -31.970 27.110 -31.720 ;
        RECT 26.860 -35.580 27.110 -35.330 ;
        RECT 26.860 -39.190 27.110 -38.940 ;
      LAYER met1 ;
        RECT 26.650 -43.100 27.330 19.120 ;
    END
  END BLb3
  PIN BL4
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER li1 ;
        RECT 28.420 14.860 28.870 15.310 ;
        RECT 28.420 11.250 28.870 11.700 ;
        RECT 28.420 7.640 28.870 8.090 ;
        RECT 28.420 4.030 28.870 4.480 ;
        RECT 28.420 0.420 28.870 0.870 ;
        RECT 28.420 -3.190 28.870 -2.740 ;
        RECT 28.420 -6.800 28.870 -6.350 ;
        RECT 28.420 -10.410 28.870 -9.960 ;
        RECT 28.420 -14.020 28.870 -13.570 ;
        RECT 28.420 -17.630 28.870 -17.180 ;
        RECT 28.420 -21.240 28.870 -20.790 ;
        RECT 28.420 -24.850 28.870 -24.400 ;
        RECT 28.420 -28.460 28.870 -28.010 ;
        RECT 28.420 -32.070 28.870 -31.620 ;
        RECT 28.420 -35.680 28.870 -35.230 ;
        RECT 28.420 -39.290 28.870 -38.840 ;
      LAYER mcon ;
        RECT 28.520 14.960 28.770 15.210 ;
        RECT 28.520 11.350 28.770 11.600 ;
        RECT 28.520 7.740 28.770 7.990 ;
        RECT 28.520 4.130 28.770 4.380 ;
        RECT 28.520 0.520 28.770 0.770 ;
        RECT 28.520 -3.090 28.770 -2.840 ;
        RECT 28.520 -6.700 28.770 -6.450 ;
        RECT 28.520 -10.310 28.770 -10.060 ;
        RECT 28.520 -13.920 28.770 -13.670 ;
        RECT 28.520 -17.530 28.770 -17.280 ;
        RECT 28.520 -21.140 28.770 -20.890 ;
        RECT 28.520 -24.750 28.770 -24.500 ;
        RECT 28.520 -28.360 28.770 -28.110 ;
        RECT 28.520 -31.970 28.770 -31.720 ;
        RECT 28.520 -35.580 28.770 -35.330 ;
        RECT 28.520 -39.190 28.770 -38.940 ;
      LAYER met1 ;
        RECT 28.300 -43.100 28.980 19.120 ;
    END
  END BL4
  PIN BLb4
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER li1 ;
        RECT 33.520 16.660 33.970 17.110 ;
        RECT 33.520 13.050 33.970 13.510 ;
        RECT 33.520 9.440 33.970 9.900 ;
        RECT 33.520 5.830 33.970 6.290 ;
        RECT 33.520 2.220 33.970 2.680 ;
        RECT 33.520 -1.390 33.970 -0.930 ;
        RECT 33.520 -5.000 33.970 -4.540 ;
        RECT 33.520 -8.610 33.970 -8.150 ;
        RECT 33.520 -12.220 33.970 -11.760 ;
        RECT 33.520 -15.830 33.970 -15.370 ;
        RECT 33.520 -19.440 33.970 -18.980 ;
        RECT 33.520 -23.050 33.970 -22.590 ;
        RECT 33.520 -26.660 33.970 -26.200 ;
        RECT 33.520 -30.270 33.970 -29.810 ;
        RECT 33.520 -33.880 33.970 -33.420 ;
        RECT 33.520 -37.490 33.970 -37.030 ;
        RECT 33.520 -41.090 33.970 -40.640 ;
      LAYER mcon ;
        RECT 33.620 16.760 33.880 17.020 ;
        RECT 33.620 13.150 33.880 13.410 ;
        RECT 33.620 9.540 33.880 9.800 ;
        RECT 33.620 5.930 33.880 6.190 ;
        RECT 33.620 2.320 33.880 2.580 ;
        RECT 33.620 -1.290 33.880 -1.030 ;
        RECT 33.620 -4.900 33.880 -4.640 ;
        RECT 33.620 -8.510 33.880 -8.250 ;
        RECT 33.620 -12.120 33.880 -11.860 ;
        RECT 33.620 -15.730 33.880 -15.470 ;
        RECT 33.620 -19.340 33.880 -19.080 ;
        RECT 33.620 -22.950 33.880 -22.690 ;
        RECT 33.620 -26.560 33.880 -26.300 ;
        RECT 33.620 -30.170 33.880 -29.910 ;
        RECT 33.620 -33.780 33.880 -33.520 ;
        RECT 33.620 -37.390 33.880 -37.130 ;
        RECT 33.620 -41.000 33.880 -40.740 ;
      LAYER met1 ;
        RECT 33.400 -43.110 34.080 19.130 ;
    END
  END BLb4
  PIN BL5
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER li1 ;
        RECT 35.160 16.660 35.610 17.110 ;
        RECT 35.160 13.050 35.610 13.510 ;
        RECT 35.160 9.440 35.610 9.900 ;
        RECT 35.160 5.830 35.610 6.290 ;
        RECT 35.160 2.220 35.610 2.680 ;
        RECT 35.160 -1.390 35.610 -0.930 ;
        RECT 35.160 -5.000 35.610 -4.540 ;
        RECT 35.160 -8.610 35.610 -8.150 ;
        RECT 35.160 -12.220 35.610 -11.760 ;
        RECT 35.160 -15.830 35.610 -15.370 ;
        RECT 35.160 -19.440 35.610 -18.980 ;
        RECT 35.160 -23.050 35.610 -22.590 ;
        RECT 35.160 -26.660 35.610 -26.200 ;
        RECT 35.160 -30.270 35.610 -29.810 ;
        RECT 35.160 -33.880 35.610 -33.420 ;
        RECT 35.160 -37.490 35.610 -37.030 ;
        RECT 35.160 -41.090 35.610 -40.640 ;
      LAYER mcon ;
        RECT 35.250 16.760 35.510 17.020 ;
        RECT 35.250 13.150 35.510 13.410 ;
        RECT 35.250 9.540 35.510 9.800 ;
        RECT 35.250 5.930 35.510 6.190 ;
        RECT 35.250 2.320 35.510 2.580 ;
        RECT 35.250 -1.290 35.510 -1.030 ;
        RECT 35.250 -4.900 35.510 -4.640 ;
        RECT 35.250 -8.510 35.510 -8.250 ;
        RECT 35.250 -12.120 35.510 -11.860 ;
        RECT 35.250 -15.730 35.510 -15.470 ;
        RECT 35.250 -19.340 35.510 -19.080 ;
        RECT 35.250 -22.950 35.510 -22.690 ;
        RECT 35.250 -26.560 35.510 -26.300 ;
        RECT 35.250 -30.170 35.510 -29.910 ;
        RECT 35.250 -33.780 35.510 -33.520 ;
        RECT 35.250 -37.390 35.510 -37.130 ;
        RECT 35.250 -41.000 35.510 -40.740 ;
      LAYER met1 ;
        RECT 35.040 -43.120 35.720 19.140 ;
    END
  END BL5
  PIN BLb5
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER li1 ;
        RECT 40.260 14.860 40.710 15.310 ;
        RECT 40.260 11.250 40.710 11.700 ;
        RECT 40.260 7.640 40.710 8.090 ;
        RECT 40.260 4.030 40.710 4.480 ;
        RECT 40.260 0.420 40.710 0.870 ;
        RECT 40.260 -3.190 40.710 -2.740 ;
        RECT 40.260 -6.800 40.710 -6.350 ;
        RECT 40.260 -10.410 40.710 -9.960 ;
        RECT 40.260 -14.020 40.710 -13.570 ;
        RECT 40.260 -17.630 40.710 -17.180 ;
        RECT 40.260 -21.240 40.710 -20.790 ;
        RECT 40.260 -24.850 40.710 -24.400 ;
        RECT 40.260 -28.460 40.710 -28.010 ;
        RECT 40.260 -32.070 40.710 -31.620 ;
        RECT 40.260 -35.680 40.710 -35.230 ;
        RECT 40.260 -39.290 40.710 -38.840 ;
      LAYER mcon ;
        RECT 40.360 14.960 40.610 15.210 ;
        RECT 40.360 11.350 40.610 11.600 ;
        RECT 40.360 7.740 40.610 7.990 ;
        RECT 40.360 4.130 40.610 4.380 ;
        RECT 40.360 0.520 40.610 0.770 ;
        RECT 40.360 -3.090 40.610 -2.840 ;
        RECT 40.360 -6.700 40.610 -6.450 ;
        RECT 40.360 -10.310 40.610 -10.060 ;
        RECT 40.360 -13.920 40.610 -13.670 ;
        RECT 40.360 -17.530 40.610 -17.280 ;
        RECT 40.360 -21.140 40.610 -20.890 ;
        RECT 40.360 -24.750 40.610 -24.500 ;
        RECT 40.360 -28.360 40.610 -28.110 ;
        RECT 40.360 -31.970 40.610 -31.720 ;
        RECT 40.360 -35.580 40.610 -35.330 ;
        RECT 40.360 -39.190 40.610 -38.940 ;
      LAYER met1 ;
        RECT 40.150 -43.110 40.830 19.130 ;
    END
  END BLb5
  PIN BL6
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER li1 ;
        RECT 41.920 14.860 42.370 15.310 ;
        RECT 41.920 11.250 42.370 11.700 ;
        RECT 41.920 7.640 42.370 8.090 ;
        RECT 41.920 4.030 42.370 4.480 ;
        RECT 41.920 0.420 42.370 0.870 ;
        RECT 41.920 -3.190 42.370 -2.740 ;
        RECT 41.920 -6.800 42.370 -6.350 ;
        RECT 41.920 -10.410 42.370 -9.960 ;
        RECT 41.920 -14.020 42.370 -13.570 ;
        RECT 41.920 -17.630 42.370 -17.180 ;
        RECT 41.920 -21.240 42.370 -20.790 ;
        RECT 41.920 -24.850 42.370 -24.400 ;
        RECT 41.920 -28.460 42.370 -28.010 ;
        RECT 41.920 -32.070 42.370 -31.620 ;
        RECT 41.920 -35.680 42.370 -35.230 ;
        RECT 41.920 -39.290 42.370 -38.840 ;
      LAYER mcon ;
        RECT 42.020 14.960 42.270 15.210 ;
        RECT 42.020 11.350 42.270 11.600 ;
        RECT 42.020 7.740 42.270 7.990 ;
        RECT 42.020 4.130 42.270 4.380 ;
        RECT 42.020 0.520 42.270 0.770 ;
        RECT 42.020 -3.090 42.270 -2.840 ;
        RECT 42.020 -6.700 42.270 -6.450 ;
        RECT 42.020 -10.310 42.270 -10.060 ;
        RECT 42.020 -13.920 42.270 -13.670 ;
        RECT 42.020 -17.530 42.270 -17.280 ;
        RECT 42.020 -21.140 42.270 -20.890 ;
        RECT 42.020 -24.750 42.270 -24.500 ;
        RECT 42.020 -28.360 42.270 -28.110 ;
        RECT 42.020 -31.970 42.270 -31.720 ;
        RECT 42.020 -35.580 42.270 -35.330 ;
        RECT 42.020 -39.190 42.270 -38.940 ;
      LAYER met1 ;
        RECT 41.790 -43.110 42.470 19.130 ;
    END
  END BL6
  PIN BLb6
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER li1 ;
        RECT 47.020 16.660 47.470 17.110 ;
        RECT 47.020 13.050 47.470 13.510 ;
        RECT 47.020 9.440 47.470 9.900 ;
        RECT 47.020 5.830 47.470 6.290 ;
        RECT 47.020 2.220 47.470 2.680 ;
        RECT 47.020 -1.390 47.470 -0.930 ;
        RECT 47.020 -5.000 47.470 -4.540 ;
        RECT 47.020 -8.610 47.470 -8.150 ;
        RECT 47.020 -12.220 47.470 -11.760 ;
        RECT 47.020 -15.830 47.470 -15.370 ;
        RECT 47.020 -19.440 47.470 -18.980 ;
        RECT 47.020 -23.050 47.470 -22.590 ;
        RECT 47.020 -26.660 47.470 -26.200 ;
        RECT 47.020 -30.270 47.470 -29.810 ;
        RECT 47.020 -33.880 47.470 -33.420 ;
        RECT 47.020 -37.490 47.470 -37.030 ;
        RECT 47.020 -41.090 47.470 -40.640 ;
      LAYER mcon ;
        RECT 47.120 16.760 47.380 17.020 ;
        RECT 47.120 13.150 47.380 13.410 ;
        RECT 47.120 9.540 47.380 9.800 ;
        RECT 47.120 5.930 47.380 6.190 ;
        RECT 47.120 2.320 47.380 2.580 ;
        RECT 47.120 -1.290 47.380 -1.030 ;
        RECT 47.120 -4.900 47.380 -4.640 ;
        RECT 47.120 -8.510 47.380 -8.250 ;
        RECT 47.120 -12.120 47.380 -11.860 ;
        RECT 47.120 -15.730 47.380 -15.470 ;
        RECT 47.120 -19.340 47.380 -19.080 ;
        RECT 47.120 -22.950 47.380 -22.690 ;
        RECT 47.120 -26.560 47.380 -26.300 ;
        RECT 47.120 -30.170 47.380 -29.910 ;
        RECT 47.120 -33.780 47.380 -33.520 ;
        RECT 47.120 -37.390 47.380 -37.130 ;
        RECT 47.120 -41.000 47.380 -40.740 ;
      LAYER met1 ;
        RECT 46.910 -43.110 47.590 19.130 ;
    END
  END BLb6
  PIN BL7
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER li1 ;
        RECT 48.660 16.660 49.110 17.110 ;
        RECT 48.660 13.050 49.110 13.510 ;
        RECT 48.660 9.440 49.110 9.900 ;
        RECT 48.660 5.830 49.110 6.290 ;
        RECT 48.660 2.220 49.110 2.680 ;
        RECT 48.660 -1.390 49.110 -0.930 ;
        RECT 48.660 -5.000 49.110 -4.540 ;
        RECT 48.660 -8.610 49.110 -8.150 ;
        RECT 48.660 -12.220 49.110 -11.760 ;
        RECT 48.660 -15.830 49.110 -15.370 ;
        RECT 48.660 -19.440 49.110 -18.980 ;
        RECT 48.660 -23.050 49.110 -22.590 ;
        RECT 48.660 -26.660 49.110 -26.200 ;
        RECT 48.660 -30.270 49.110 -29.810 ;
        RECT 48.660 -33.880 49.110 -33.420 ;
        RECT 48.660 -37.490 49.110 -37.030 ;
        RECT 48.660 -41.090 49.110 -40.640 ;
      LAYER mcon ;
        RECT 48.750 16.760 49.010 17.020 ;
        RECT 48.750 13.150 49.010 13.410 ;
        RECT 48.750 9.540 49.010 9.800 ;
        RECT 48.750 5.930 49.010 6.190 ;
        RECT 48.750 2.320 49.010 2.580 ;
        RECT 48.750 -1.290 49.010 -1.030 ;
        RECT 48.750 -4.900 49.010 -4.640 ;
        RECT 48.750 -8.510 49.010 -8.250 ;
        RECT 48.750 -12.120 49.010 -11.860 ;
        RECT 48.750 -15.730 49.010 -15.470 ;
        RECT 48.750 -19.340 49.010 -19.080 ;
        RECT 48.750 -22.950 49.010 -22.690 ;
        RECT 48.750 -26.560 49.010 -26.300 ;
        RECT 48.750 -30.170 49.010 -29.910 ;
        RECT 48.750 -33.780 49.010 -33.520 ;
        RECT 48.750 -37.390 49.010 -37.130 ;
        RECT 48.750 -41.000 49.010 -40.740 ;
      LAYER met1 ;
        RECT 48.550 -43.120 49.230 19.140 ;
    END
  END BL7
  PIN BLb7
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER li1 ;
        RECT 53.760 14.860 54.210 15.310 ;
        RECT 53.760 11.250 54.210 11.700 ;
        RECT 53.760 7.640 54.210 8.090 ;
        RECT 53.760 4.030 54.210 4.480 ;
        RECT 53.760 0.420 54.210 0.870 ;
        RECT 53.760 -3.190 54.210 -2.740 ;
        RECT 53.760 -6.800 54.210 -6.350 ;
        RECT 53.760 -10.410 54.210 -9.960 ;
        RECT 53.760 -14.020 54.210 -13.570 ;
        RECT 53.760 -17.630 54.210 -17.180 ;
        RECT 53.760 -21.240 54.210 -20.790 ;
        RECT 53.760 -24.850 54.210 -24.400 ;
        RECT 53.760 -28.460 54.210 -28.010 ;
        RECT 53.760 -32.070 54.210 -31.620 ;
        RECT 53.760 -35.680 54.210 -35.230 ;
        RECT 53.760 -39.290 54.210 -38.840 ;
      LAYER mcon ;
        RECT 53.860 14.960 54.110 15.210 ;
        RECT 53.860 11.350 54.110 11.600 ;
        RECT 53.860 7.740 54.110 7.990 ;
        RECT 53.860 4.130 54.110 4.380 ;
        RECT 53.860 0.520 54.110 0.770 ;
        RECT 53.860 -3.090 54.110 -2.840 ;
        RECT 53.860 -6.700 54.110 -6.450 ;
        RECT 53.860 -10.310 54.110 -10.060 ;
        RECT 53.860 -13.920 54.110 -13.670 ;
        RECT 53.860 -17.530 54.110 -17.280 ;
        RECT 53.860 -21.140 54.110 -20.890 ;
        RECT 53.860 -24.750 54.110 -24.500 ;
        RECT 53.860 -28.360 54.110 -28.110 ;
        RECT 53.860 -31.970 54.110 -31.720 ;
        RECT 53.860 -35.580 54.110 -35.330 ;
        RECT 53.860 -39.190 54.110 -38.940 ;
      LAYER met1 ;
        RECT 53.650 -43.100 54.330 19.120 ;
    END
  END BLb7
  PIN BL8
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER li1 ;
        RECT 55.420 14.860 55.870 15.310 ;
        RECT 55.420 11.250 55.870 11.700 ;
        RECT 55.420 7.640 55.870 8.090 ;
        RECT 55.420 4.030 55.870 4.480 ;
        RECT 55.420 0.420 55.870 0.870 ;
        RECT 55.420 -3.190 55.870 -2.740 ;
        RECT 55.420 -6.800 55.870 -6.350 ;
        RECT 55.420 -10.410 55.870 -9.960 ;
        RECT 55.420 -14.020 55.870 -13.570 ;
        RECT 55.420 -17.630 55.870 -17.180 ;
        RECT 55.420 -21.240 55.870 -20.790 ;
        RECT 55.420 -24.850 55.870 -24.400 ;
        RECT 55.420 -28.460 55.870 -28.010 ;
        RECT 55.420 -32.070 55.870 -31.620 ;
        RECT 55.420 -35.680 55.870 -35.230 ;
        RECT 55.420 -39.290 55.870 -38.840 ;
      LAYER mcon ;
        RECT 55.520 14.960 55.770 15.210 ;
        RECT 55.520 11.350 55.770 11.600 ;
        RECT 55.520 7.740 55.770 7.990 ;
        RECT 55.520 4.130 55.770 4.380 ;
        RECT 55.520 0.520 55.770 0.770 ;
        RECT 55.520 -3.090 55.770 -2.840 ;
        RECT 55.520 -6.700 55.770 -6.450 ;
        RECT 55.520 -10.310 55.770 -10.060 ;
        RECT 55.520 -13.920 55.770 -13.670 ;
        RECT 55.520 -17.530 55.770 -17.280 ;
        RECT 55.520 -21.140 55.770 -20.890 ;
        RECT 55.520 -24.750 55.770 -24.500 ;
        RECT 55.520 -28.360 55.770 -28.110 ;
        RECT 55.520 -31.970 55.770 -31.720 ;
        RECT 55.520 -35.580 55.770 -35.330 ;
        RECT 55.520 -39.190 55.770 -38.940 ;
      LAYER met1 ;
        RECT 55.300 -43.100 55.980 19.120 ;
    END
  END BL8
  PIN BLb8
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER li1 ;
        RECT 60.520 16.660 60.970 17.110 ;
        RECT 60.520 13.050 60.970 13.510 ;
        RECT 60.520 9.440 60.970 9.900 ;
        RECT 60.520 5.830 60.970 6.290 ;
        RECT 60.520 2.220 60.970 2.680 ;
        RECT 60.520 -1.390 60.970 -0.930 ;
        RECT 60.520 -5.000 60.970 -4.540 ;
        RECT 60.520 -8.610 60.970 -8.150 ;
        RECT 60.520 -12.220 60.970 -11.760 ;
        RECT 60.520 -15.830 60.970 -15.370 ;
        RECT 60.520 -19.440 60.970 -18.980 ;
        RECT 60.520 -23.050 60.970 -22.590 ;
        RECT 60.520 -26.660 60.970 -26.200 ;
        RECT 60.520 -30.270 60.970 -29.810 ;
        RECT 60.520 -33.880 60.970 -33.420 ;
        RECT 60.520 -37.490 60.970 -37.030 ;
        RECT 60.520 -41.090 60.970 -40.640 ;
      LAYER mcon ;
        RECT 60.620 16.760 60.880 17.020 ;
        RECT 60.620 13.150 60.880 13.410 ;
        RECT 60.620 9.540 60.880 9.800 ;
        RECT 60.620 5.930 60.880 6.190 ;
        RECT 60.620 2.320 60.880 2.580 ;
        RECT 60.620 -1.290 60.880 -1.030 ;
        RECT 60.620 -4.900 60.880 -4.640 ;
        RECT 60.620 -8.510 60.880 -8.250 ;
        RECT 60.620 -12.120 60.880 -11.860 ;
        RECT 60.620 -15.730 60.880 -15.470 ;
        RECT 60.620 -19.340 60.880 -19.080 ;
        RECT 60.620 -22.950 60.880 -22.690 ;
        RECT 60.620 -26.560 60.880 -26.300 ;
        RECT 60.620 -30.170 60.880 -29.910 ;
        RECT 60.620 -33.780 60.880 -33.520 ;
        RECT 60.620 -37.390 60.880 -37.130 ;
        RECT 60.620 -41.000 60.880 -40.740 ;
      LAYER met1 ;
        RECT 60.400 -43.120 61.080 19.140 ;
    END
  END BLb8
  PIN BL9
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER li1 ;
        RECT 62.160 16.660 62.610 17.110 ;
        RECT 62.160 13.050 62.610 13.510 ;
        RECT 62.160 9.440 62.610 9.900 ;
        RECT 62.160 5.830 62.610 6.290 ;
        RECT 62.160 2.220 62.610 2.680 ;
        RECT 62.160 -1.390 62.610 -0.930 ;
        RECT 62.160 -5.000 62.610 -4.540 ;
        RECT 62.160 -8.610 62.610 -8.150 ;
        RECT 62.160 -12.220 62.610 -11.760 ;
        RECT 62.160 -15.830 62.610 -15.370 ;
        RECT 62.160 -19.440 62.610 -18.980 ;
        RECT 62.160 -23.050 62.610 -22.590 ;
        RECT 62.160 -26.660 62.610 -26.200 ;
        RECT 62.160 -30.270 62.610 -29.810 ;
        RECT 62.160 -33.880 62.610 -33.420 ;
        RECT 62.160 -37.490 62.610 -37.030 ;
        RECT 62.160 -41.090 62.610 -40.640 ;
      LAYER mcon ;
        RECT 62.250 16.760 62.510 17.020 ;
        RECT 62.250 13.150 62.510 13.410 ;
        RECT 62.250 9.540 62.510 9.800 ;
        RECT 62.250 5.930 62.510 6.190 ;
        RECT 62.250 2.320 62.510 2.580 ;
        RECT 62.250 -1.290 62.510 -1.030 ;
        RECT 62.250 -4.900 62.510 -4.640 ;
        RECT 62.250 -8.510 62.510 -8.250 ;
        RECT 62.250 -12.120 62.510 -11.860 ;
        RECT 62.250 -15.730 62.510 -15.470 ;
        RECT 62.250 -19.340 62.510 -19.080 ;
        RECT 62.250 -22.950 62.510 -22.690 ;
        RECT 62.250 -26.560 62.510 -26.300 ;
        RECT 62.250 -30.170 62.510 -29.910 ;
        RECT 62.250 -33.780 62.510 -33.520 ;
        RECT 62.250 -37.390 62.510 -37.130 ;
        RECT 62.250 -41.000 62.510 -40.740 ;
      LAYER met1 ;
        RECT 62.040 -43.110 62.720 19.130 ;
    END
  END BL9
  PIN BLb9
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER li1 ;
        RECT 67.260 14.860 67.710 15.310 ;
        RECT 67.260 11.250 67.710 11.700 ;
        RECT 67.260 7.640 67.710 8.090 ;
        RECT 67.260 4.030 67.710 4.480 ;
        RECT 67.260 0.420 67.710 0.870 ;
        RECT 67.260 -3.190 67.710 -2.740 ;
        RECT 67.260 -6.800 67.710 -6.350 ;
        RECT 67.260 -10.410 67.710 -9.960 ;
        RECT 67.260 -14.020 67.710 -13.570 ;
        RECT 67.260 -17.630 67.710 -17.180 ;
        RECT 67.260 -21.240 67.710 -20.790 ;
        RECT 67.260 -24.850 67.710 -24.400 ;
        RECT 67.260 -28.460 67.710 -28.010 ;
        RECT 67.260 -32.070 67.710 -31.620 ;
        RECT 67.260 -35.680 67.710 -35.230 ;
        RECT 67.260 -39.290 67.710 -38.840 ;
      LAYER mcon ;
        RECT 67.360 14.960 67.610 15.210 ;
        RECT 67.360 11.350 67.610 11.600 ;
        RECT 67.360 7.740 67.610 7.990 ;
        RECT 67.360 4.130 67.610 4.380 ;
        RECT 67.360 0.520 67.610 0.770 ;
        RECT 67.360 -3.090 67.610 -2.840 ;
        RECT 67.360 -6.700 67.610 -6.450 ;
        RECT 67.360 -10.310 67.610 -10.060 ;
        RECT 67.360 -13.920 67.610 -13.670 ;
        RECT 67.360 -17.530 67.610 -17.280 ;
        RECT 67.360 -21.140 67.610 -20.890 ;
        RECT 67.360 -24.750 67.610 -24.500 ;
        RECT 67.360 -28.360 67.610 -28.110 ;
        RECT 67.360 -31.970 67.610 -31.720 ;
        RECT 67.360 -35.580 67.610 -35.330 ;
        RECT 67.360 -39.190 67.610 -38.940 ;
      LAYER met1 ;
        RECT 67.330 19.130 67.680 19.140 ;
        RECT 67.160 -43.110 67.840 19.130 ;
    END
  END BLb9
  PIN BL10
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER li1 ;
        RECT 68.920 14.860 69.370 15.310 ;
        RECT 68.920 11.250 69.370 11.700 ;
        RECT 68.920 7.640 69.370 8.090 ;
        RECT 68.920 4.030 69.370 4.480 ;
        RECT 68.920 0.420 69.370 0.870 ;
        RECT 68.920 -3.190 69.370 -2.740 ;
        RECT 68.920 -6.800 69.370 -6.350 ;
        RECT 68.920 -10.410 69.370 -9.960 ;
        RECT 68.920 -14.020 69.370 -13.570 ;
        RECT 68.920 -17.630 69.370 -17.180 ;
        RECT 68.920 -21.240 69.370 -20.790 ;
        RECT 68.920 -24.850 69.370 -24.400 ;
        RECT 68.920 -28.460 69.370 -28.010 ;
        RECT 68.920 -32.070 69.370 -31.620 ;
        RECT 68.920 -35.680 69.370 -35.230 ;
        RECT 68.920 -39.290 69.370 -38.840 ;
      LAYER mcon ;
        RECT 69.020 14.960 69.270 15.210 ;
        RECT 69.020 11.350 69.270 11.600 ;
        RECT 69.020 7.740 69.270 7.990 ;
        RECT 69.020 4.130 69.270 4.380 ;
        RECT 69.020 0.520 69.270 0.770 ;
        RECT 69.020 -3.090 69.270 -2.840 ;
        RECT 69.020 -6.700 69.270 -6.450 ;
        RECT 69.020 -10.310 69.270 -10.060 ;
        RECT 69.020 -13.920 69.270 -13.670 ;
        RECT 69.020 -17.530 69.270 -17.280 ;
        RECT 69.020 -21.140 69.270 -20.890 ;
        RECT 69.020 -24.750 69.270 -24.500 ;
        RECT 69.020 -28.360 69.270 -28.110 ;
        RECT 69.020 -31.970 69.270 -31.720 ;
        RECT 69.020 -35.580 69.270 -35.330 ;
        RECT 69.020 -39.190 69.270 -38.940 ;
      LAYER met1 ;
        RECT 68.800 -43.110 69.480 19.130 ;
    END
  END BL10
  PIN BLb10
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER li1 ;
        RECT 74.020 16.660 74.470 17.110 ;
        RECT 74.020 13.050 74.470 13.510 ;
        RECT 74.020 9.440 74.470 9.900 ;
        RECT 74.020 5.830 74.470 6.290 ;
        RECT 74.020 2.220 74.470 2.680 ;
        RECT 74.020 -1.390 74.470 -0.930 ;
        RECT 74.020 -5.000 74.470 -4.540 ;
        RECT 74.020 -8.610 74.470 -8.150 ;
        RECT 74.020 -12.220 74.470 -11.760 ;
        RECT 74.020 -15.830 74.470 -15.370 ;
        RECT 74.020 -19.440 74.470 -18.980 ;
        RECT 74.020 -23.050 74.470 -22.590 ;
        RECT 74.020 -26.660 74.470 -26.200 ;
        RECT 74.020 -30.270 74.470 -29.810 ;
        RECT 74.020 -33.880 74.470 -33.420 ;
        RECT 74.020 -37.490 74.470 -37.030 ;
        RECT 74.020 -41.090 74.470 -40.640 ;
      LAYER mcon ;
        RECT 74.120 16.760 74.380 17.020 ;
        RECT 74.120 13.150 74.380 13.410 ;
        RECT 74.120 9.540 74.380 9.800 ;
        RECT 74.120 5.930 74.380 6.190 ;
        RECT 74.120 2.320 74.380 2.580 ;
        RECT 74.120 -1.290 74.380 -1.030 ;
        RECT 74.120 -4.900 74.380 -4.640 ;
        RECT 74.120 -8.510 74.380 -8.250 ;
        RECT 74.120 -12.120 74.380 -11.860 ;
        RECT 74.120 -15.730 74.380 -15.470 ;
        RECT 74.120 -19.340 74.380 -19.080 ;
        RECT 74.120 -22.950 74.380 -22.690 ;
        RECT 74.120 -26.560 74.380 -26.300 ;
        RECT 74.120 -30.170 74.380 -29.910 ;
        RECT 74.120 -33.780 74.380 -33.520 ;
        RECT 74.120 -37.390 74.380 -37.130 ;
        RECT 74.120 -41.000 74.380 -40.740 ;
      LAYER met1 ;
        RECT 73.910 -43.120 74.590 19.140 ;
    END
  END BLb10
  PIN BL11
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER li1 ;
        RECT 75.660 16.660 76.110 17.110 ;
        RECT 75.660 13.050 76.110 13.510 ;
        RECT 75.660 9.440 76.110 9.900 ;
        RECT 75.660 5.830 76.110 6.290 ;
        RECT 75.660 2.220 76.110 2.680 ;
        RECT 75.660 -1.390 76.110 -0.930 ;
        RECT 75.660 -5.000 76.110 -4.540 ;
        RECT 75.660 -8.610 76.110 -8.150 ;
        RECT 75.660 -12.220 76.110 -11.760 ;
        RECT 75.660 -15.830 76.110 -15.370 ;
        RECT 75.660 -19.440 76.110 -18.980 ;
        RECT 75.660 -23.050 76.110 -22.590 ;
        RECT 75.660 -26.660 76.110 -26.200 ;
        RECT 75.660 -30.270 76.110 -29.810 ;
        RECT 75.660 -33.880 76.110 -33.420 ;
        RECT 75.660 -37.490 76.110 -37.030 ;
        RECT 75.660 -41.090 76.110 -40.640 ;
      LAYER mcon ;
        RECT 75.750 16.760 76.010 17.020 ;
        RECT 75.750 13.150 76.010 13.410 ;
        RECT 75.750 9.540 76.010 9.800 ;
        RECT 75.750 5.930 76.010 6.190 ;
        RECT 75.750 2.320 76.010 2.580 ;
        RECT 75.750 -1.290 76.010 -1.030 ;
        RECT 75.750 -4.900 76.010 -4.640 ;
        RECT 75.750 -8.510 76.010 -8.250 ;
        RECT 75.750 -12.120 76.010 -11.860 ;
        RECT 75.750 -15.730 76.010 -15.470 ;
        RECT 75.750 -19.340 76.010 -19.080 ;
        RECT 75.750 -22.950 76.010 -22.690 ;
        RECT 75.750 -26.560 76.010 -26.300 ;
        RECT 75.750 -30.170 76.010 -29.910 ;
        RECT 75.750 -33.780 76.010 -33.520 ;
        RECT 75.750 -37.390 76.010 -37.130 ;
        RECT 75.750 -41.000 76.010 -40.740 ;
      LAYER met1 ;
        RECT 75.550 -43.110 76.230 19.130 ;
    END
  END BL11
  PIN BLb11
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER li1 ;
        RECT 80.760 14.860 81.210 15.310 ;
        RECT 80.760 11.250 81.210 11.700 ;
        RECT 80.760 7.640 81.210 8.090 ;
        RECT 80.760 4.030 81.210 4.480 ;
        RECT 80.760 0.420 81.210 0.870 ;
        RECT 80.760 -3.190 81.210 -2.740 ;
        RECT 80.760 -6.800 81.210 -6.350 ;
        RECT 80.760 -10.410 81.210 -9.960 ;
        RECT 80.760 -14.020 81.210 -13.570 ;
        RECT 80.760 -17.630 81.210 -17.180 ;
        RECT 80.760 -21.240 81.210 -20.790 ;
        RECT 80.760 -24.850 81.210 -24.400 ;
        RECT 80.760 -28.460 81.210 -28.010 ;
        RECT 80.760 -32.070 81.210 -31.620 ;
        RECT 80.760 -35.680 81.210 -35.230 ;
        RECT 80.760 -39.290 81.210 -38.840 ;
      LAYER mcon ;
        RECT 80.860 14.960 81.110 15.210 ;
        RECT 80.860 11.350 81.110 11.600 ;
        RECT 80.860 7.740 81.110 7.990 ;
        RECT 80.860 4.130 81.110 4.380 ;
        RECT 80.860 0.520 81.110 0.770 ;
        RECT 80.860 -3.090 81.110 -2.840 ;
        RECT 80.860 -6.700 81.110 -6.450 ;
        RECT 80.860 -10.310 81.110 -10.060 ;
        RECT 80.860 -13.920 81.110 -13.670 ;
        RECT 80.860 -17.530 81.110 -17.280 ;
        RECT 80.860 -21.140 81.110 -20.890 ;
        RECT 80.860 -24.750 81.110 -24.500 ;
        RECT 80.860 -28.360 81.110 -28.110 ;
        RECT 80.860 -31.970 81.110 -31.720 ;
        RECT 80.860 -35.580 81.110 -35.330 ;
        RECT 80.860 -39.190 81.110 -38.940 ;
      LAYER met1 ;
        RECT 80.830 19.120 81.180 19.130 ;
        RECT 80.650 -43.100 81.330 19.120 ;
    END
  END BLb11
  PIN BL12
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER li1 ;
        RECT 82.420 14.860 82.870 15.310 ;
        RECT 82.420 11.250 82.870 11.700 ;
        RECT 82.420 7.640 82.870 8.090 ;
        RECT 82.420 4.030 82.870 4.480 ;
        RECT 82.420 0.420 82.870 0.870 ;
        RECT 82.420 -3.190 82.870 -2.740 ;
        RECT 82.420 -6.800 82.870 -6.350 ;
        RECT 82.420 -10.410 82.870 -9.960 ;
        RECT 82.420 -14.020 82.870 -13.570 ;
        RECT 82.420 -17.630 82.870 -17.180 ;
        RECT 82.420 -21.240 82.870 -20.790 ;
        RECT 82.420 -24.850 82.870 -24.400 ;
        RECT 82.420 -28.460 82.870 -28.010 ;
        RECT 82.420 -32.070 82.870 -31.620 ;
        RECT 82.420 -35.680 82.870 -35.230 ;
        RECT 82.420 -39.290 82.870 -38.840 ;
      LAYER mcon ;
        RECT 82.520 14.960 82.770 15.210 ;
        RECT 82.520 11.350 82.770 11.600 ;
        RECT 82.520 7.740 82.770 7.990 ;
        RECT 82.520 4.130 82.770 4.380 ;
        RECT 82.520 0.520 82.770 0.770 ;
        RECT 82.520 -3.090 82.770 -2.840 ;
        RECT 82.520 -6.700 82.770 -6.450 ;
        RECT 82.520 -10.310 82.770 -10.060 ;
        RECT 82.520 -13.920 82.770 -13.670 ;
        RECT 82.520 -17.530 82.770 -17.280 ;
        RECT 82.520 -21.140 82.770 -20.890 ;
        RECT 82.520 -24.750 82.770 -24.500 ;
        RECT 82.520 -28.360 82.770 -28.110 ;
        RECT 82.520 -31.970 82.770 -31.720 ;
        RECT 82.520 -35.580 82.770 -35.330 ;
        RECT 82.520 -39.190 82.770 -38.940 ;
      LAYER met1 ;
        RECT 82.300 -43.100 82.980 19.120 ;
    END
  END BL12
  PIN BLb12
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER li1 ;
        RECT 87.520 16.660 87.970 17.110 ;
        RECT 87.520 13.050 87.970 13.510 ;
        RECT 87.520 9.440 87.970 9.900 ;
        RECT 87.520 5.830 87.970 6.290 ;
        RECT 87.520 2.220 87.970 2.680 ;
        RECT 87.520 -1.390 87.970 -0.930 ;
        RECT 87.520 -5.000 87.970 -4.540 ;
        RECT 87.520 -8.610 87.970 -8.150 ;
        RECT 87.520 -12.220 87.970 -11.760 ;
        RECT 87.520 -15.830 87.970 -15.370 ;
        RECT 87.520 -19.440 87.970 -18.980 ;
        RECT 87.520 -23.050 87.970 -22.590 ;
        RECT 87.520 -26.660 87.970 -26.200 ;
        RECT 87.520 -30.270 87.970 -29.810 ;
        RECT 87.520 -33.880 87.970 -33.420 ;
        RECT 87.520 -37.490 87.970 -37.030 ;
        RECT 87.520 -41.090 87.970 -40.640 ;
      LAYER mcon ;
        RECT 87.620 16.760 87.880 17.020 ;
        RECT 87.620 13.150 87.880 13.410 ;
        RECT 87.620 9.540 87.880 9.800 ;
        RECT 87.620 5.930 87.880 6.190 ;
        RECT 87.620 2.320 87.880 2.580 ;
        RECT 87.620 -1.290 87.880 -1.030 ;
        RECT 87.620 -4.900 87.880 -4.640 ;
        RECT 87.620 -8.510 87.880 -8.250 ;
        RECT 87.620 -12.120 87.880 -11.860 ;
        RECT 87.620 -15.730 87.880 -15.470 ;
        RECT 87.620 -19.340 87.880 -19.080 ;
        RECT 87.620 -22.950 87.880 -22.690 ;
        RECT 87.620 -26.560 87.880 -26.300 ;
        RECT 87.620 -30.170 87.880 -29.910 ;
        RECT 87.620 -33.780 87.880 -33.520 ;
        RECT 87.620 -37.390 87.880 -37.130 ;
        RECT 87.620 -41.000 87.880 -40.740 ;
      LAYER met1 ;
        RECT 87.400 -43.110 88.080 19.130 ;
    END
  END BLb12
  PIN BL13
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER li1 ;
        RECT 89.160 16.660 89.610 17.110 ;
        RECT 89.160 13.050 89.610 13.510 ;
        RECT 89.160 9.440 89.610 9.900 ;
        RECT 89.160 5.830 89.610 6.290 ;
        RECT 89.160 2.220 89.610 2.680 ;
        RECT 89.160 -1.390 89.610 -0.930 ;
        RECT 89.160 -5.000 89.610 -4.540 ;
        RECT 89.160 -8.610 89.610 -8.150 ;
        RECT 89.160 -12.220 89.610 -11.760 ;
        RECT 89.160 -15.830 89.610 -15.370 ;
        RECT 89.160 -19.440 89.610 -18.980 ;
        RECT 89.160 -23.050 89.610 -22.590 ;
        RECT 89.160 -26.660 89.610 -26.200 ;
        RECT 89.160 -30.270 89.610 -29.810 ;
        RECT 89.160 -33.880 89.610 -33.420 ;
        RECT 89.160 -37.490 89.610 -37.030 ;
        RECT 89.160 -41.090 89.610 -40.640 ;
      LAYER mcon ;
        RECT 89.250 16.760 89.510 17.020 ;
        RECT 89.250 13.150 89.510 13.410 ;
        RECT 89.250 9.540 89.510 9.800 ;
        RECT 89.250 5.930 89.510 6.190 ;
        RECT 89.250 2.320 89.510 2.580 ;
        RECT 89.250 -1.290 89.510 -1.030 ;
        RECT 89.250 -4.900 89.510 -4.640 ;
        RECT 89.250 -8.510 89.510 -8.250 ;
        RECT 89.250 -12.120 89.510 -11.860 ;
        RECT 89.250 -15.730 89.510 -15.470 ;
        RECT 89.250 -19.340 89.510 -19.080 ;
        RECT 89.250 -22.950 89.510 -22.690 ;
        RECT 89.250 -26.560 89.510 -26.300 ;
        RECT 89.250 -30.170 89.510 -29.910 ;
        RECT 89.250 -33.780 89.510 -33.520 ;
        RECT 89.250 -37.390 89.510 -37.130 ;
        RECT 89.250 -41.000 89.510 -40.740 ;
      LAYER met1 ;
        RECT 89.040 -43.120 89.720 19.140 ;
    END
  END BL13
  PIN BLb13
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER li1 ;
        RECT 94.260 14.860 94.710 15.310 ;
        RECT 94.260 11.250 94.710 11.700 ;
        RECT 94.260 7.640 94.710 8.090 ;
        RECT 94.260 4.030 94.710 4.480 ;
        RECT 94.260 0.420 94.710 0.870 ;
        RECT 94.260 -3.190 94.710 -2.740 ;
        RECT 94.260 -6.800 94.710 -6.350 ;
        RECT 94.260 -10.410 94.710 -9.960 ;
        RECT 94.260 -14.020 94.710 -13.570 ;
        RECT 94.260 -17.630 94.710 -17.180 ;
        RECT 94.260 -21.240 94.710 -20.790 ;
        RECT 94.260 -24.850 94.710 -24.400 ;
        RECT 94.260 -28.460 94.710 -28.010 ;
        RECT 94.260 -32.070 94.710 -31.620 ;
        RECT 94.260 -35.680 94.710 -35.230 ;
        RECT 94.260 -39.290 94.710 -38.840 ;
      LAYER mcon ;
        RECT 94.360 14.960 94.610 15.210 ;
        RECT 94.360 11.350 94.610 11.600 ;
        RECT 94.360 7.740 94.610 7.990 ;
        RECT 94.360 4.130 94.610 4.380 ;
        RECT 94.360 0.520 94.610 0.770 ;
        RECT 94.360 -3.090 94.610 -2.840 ;
        RECT 94.360 -6.700 94.610 -6.450 ;
        RECT 94.360 -10.310 94.610 -10.060 ;
        RECT 94.360 -13.920 94.610 -13.670 ;
        RECT 94.360 -17.530 94.610 -17.280 ;
        RECT 94.360 -21.140 94.610 -20.890 ;
        RECT 94.360 -24.750 94.610 -24.500 ;
        RECT 94.360 -28.360 94.610 -28.110 ;
        RECT 94.360 -31.970 94.610 -31.720 ;
        RECT 94.360 -35.580 94.610 -35.330 ;
        RECT 94.360 -39.190 94.610 -38.940 ;
      LAYER met1 ;
        RECT 94.150 -43.110 94.830 19.130 ;
    END
  END BLb13
  PIN BL14
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER li1 ;
        RECT 95.920 14.860 96.370 15.310 ;
        RECT 95.920 11.250 96.370 11.700 ;
        RECT 95.920 7.640 96.370 8.090 ;
        RECT 95.920 4.030 96.370 4.480 ;
        RECT 95.920 0.420 96.370 0.870 ;
        RECT 95.920 -3.190 96.370 -2.740 ;
        RECT 95.920 -6.800 96.370 -6.350 ;
        RECT 95.920 -10.410 96.370 -9.960 ;
        RECT 95.920 -14.020 96.370 -13.570 ;
        RECT 95.920 -17.630 96.370 -17.180 ;
        RECT 95.920 -21.240 96.370 -20.790 ;
        RECT 95.920 -24.850 96.370 -24.400 ;
        RECT 95.920 -28.460 96.370 -28.010 ;
        RECT 95.920 -32.070 96.370 -31.620 ;
        RECT 95.920 -35.680 96.370 -35.230 ;
        RECT 95.920 -39.290 96.370 -38.840 ;
      LAYER mcon ;
        RECT 96.020 14.960 96.270 15.210 ;
        RECT 96.020 11.350 96.270 11.600 ;
        RECT 96.020 7.740 96.270 7.990 ;
        RECT 96.020 4.130 96.270 4.380 ;
        RECT 96.020 0.520 96.270 0.770 ;
        RECT 96.020 -3.090 96.270 -2.840 ;
        RECT 96.020 -6.700 96.270 -6.450 ;
        RECT 96.020 -10.310 96.270 -10.060 ;
        RECT 96.020 -13.920 96.270 -13.670 ;
        RECT 96.020 -17.530 96.270 -17.280 ;
        RECT 96.020 -21.140 96.270 -20.890 ;
        RECT 96.020 -24.750 96.270 -24.500 ;
        RECT 96.020 -28.360 96.270 -28.110 ;
        RECT 96.020 -31.970 96.270 -31.720 ;
        RECT 96.020 -35.580 96.270 -35.330 ;
        RECT 96.020 -39.190 96.270 -38.940 ;
      LAYER met1 ;
        RECT 95.790 -43.110 96.470 19.130 ;
    END
  END BL14
  PIN BLb14
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER li1 ;
        RECT 101.020 16.660 101.470 17.110 ;
        RECT 101.020 13.050 101.470 13.510 ;
        RECT 101.020 9.440 101.470 9.900 ;
        RECT 101.020 5.830 101.470 6.290 ;
        RECT 101.020 2.220 101.470 2.680 ;
        RECT 101.020 -1.390 101.470 -0.930 ;
        RECT 101.020 -5.000 101.470 -4.540 ;
        RECT 101.020 -8.610 101.470 -8.150 ;
        RECT 101.020 -12.220 101.470 -11.760 ;
        RECT 101.020 -15.830 101.470 -15.370 ;
        RECT 101.020 -19.440 101.470 -18.980 ;
        RECT 101.020 -23.050 101.470 -22.590 ;
        RECT 101.020 -26.660 101.470 -26.200 ;
        RECT 101.020 -30.270 101.470 -29.810 ;
        RECT 101.020 -33.880 101.470 -33.420 ;
        RECT 101.020 -37.490 101.470 -37.030 ;
        RECT 101.020 -41.090 101.470 -40.640 ;
      LAYER mcon ;
        RECT 101.120 16.760 101.380 17.020 ;
        RECT 101.120 13.150 101.380 13.410 ;
        RECT 101.120 9.540 101.380 9.800 ;
        RECT 101.120 5.930 101.380 6.190 ;
        RECT 101.120 2.320 101.380 2.580 ;
        RECT 101.120 -1.290 101.380 -1.030 ;
        RECT 101.120 -4.900 101.380 -4.640 ;
        RECT 101.120 -8.510 101.380 -8.250 ;
        RECT 101.120 -12.120 101.380 -11.860 ;
        RECT 101.120 -15.730 101.380 -15.470 ;
        RECT 101.120 -19.340 101.380 -19.080 ;
        RECT 101.120 -22.950 101.380 -22.690 ;
        RECT 101.120 -26.560 101.380 -26.300 ;
        RECT 101.120 -30.170 101.380 -29.910 ;
        RECT 101.120 -33.780 101.380 -33.520 ;
        RECT 101.120 -37.390 101.380 -37.130 ;
        RECT 101.120 -41.000 101.380 -40.740 ;
      LAYER met1 ;
        RECT 100.910 -43.110 101.590 19.130 ;
    END
  END BLb14
  PIN BL15
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER li1 ;
        RECT 102.660 16.660 103.110 17.110 ;
        RECT 102.660 13.050 103.110 13.510 ;
        RECT 102.660 9.440 103.110 9.900 ;
        RECT 102.660 5.830 103.110 6.290 ;
        RECT 102.660 2.220 103.110 2.680 ;
        RECT 102.660 -1.390 103.110 -0.930 ;
        RECT 102.660 -5.000 103.110 -4.540 ;
        RECT 102.660 -8.610 103.110 -8.150 ;
        RECT 102.660 -12.220 103.110 -11.760 ;
        RECT 102.660 -15.830 103.110 -15.370 ;
        RECT 102.660 -19.440 103.110 -18.980 ;
        RECT 102.660 -23.050 103.110 -22.590 ;
        RECT 102.660 -26.660 103.110 -26.200 ;
        RECT 102.660 -30.270 103.110 -29.810 ;
        RECT 102.660 -33.880 103.110 -33.420 ;
        RECT 102.660 -37.490 103.110 -37.030 ;
        RECT 102.660 -41.090 103.110 -40.640 ;
      LAYER mcon ;
        RECT 102.750 16.760 103.010 17.020 ;
        RECT 102.750 13.150 103.010 13.410 ;
        RECT 102.750 9.540 103.010 9.800 ;
        RECT 102.750 5.930 103.010 6.190 ;
        RECT 102.750 2.320 103.010 2.580 ;
        RECT 102.750 -1.290 103.010 -1.030 ;
        RECT 102.750 -4.900 103.010 -4.640 ;
        RECT 102.750 -8.510 103.010 -8.250 ;
        RECT 102.750 -12.120 103.010 -11.860 ;
        RECT 102.750 -15.730 103.010 -15.470 ;
        RECT 102.750 -19.340 103.010 -19.080 ;
        RECT 102.750 -22.950 103.010 -22.690 ;
        RECT 102.750 -26.560 103.010 -26.300 ;
        RECT 102.750 -30.170 103.010 -29.910 ;
        RECT 102.750 -33.780 103.010 -33.520 ;
        RECT 102.750 -37.390 103.010 -37.130 ;
        RECT 102.750 -41.000 103.010 -40.740 ;
      LAYER met1 ;
        RECT 102.550 -43.120 103.230 19.140 ;
    END
  END BL15
  PIN BLb15
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER li1 ;
        RECT 107.760 14.860 108.210 15.310 ;
        RECT 107.760 11.250 108.210 11.700 ;
        RECT 107.760 7.640 108.210 8.090 ;
        RECT 107.760 4.030 108.210 4.480 ;
        RECT 107.760 0.420 108.210 0.870 ;
        RECT 107.760 -3.190 108.210 -2.740 ;
        RECT 107.760 -6.800 108.210 -6.350 ;
        RECT 107.760 -10.410 108.210 -9.960 ;
        RECT 107.760 -14.020 108.210 -13.570 ;
        RECT 107.760 -17.630 108.210 -17.180 ;
        RECT 107.760 -21.240 108.210 -20.790 ;
        RECT 107.760 -24.850 108.210 -24.400 ;
        RECT 107.760 -28.460 108.210 -28.010 ;
        RECT 107.760 -32.070 108.210 -31.620 ;
        RECT 107.760 -35.680 108.210 -35.230 ;
        RECT 107.760 -39.290 108.210 -38.840 ;
      LAYER mcon ;
        RECT 107.860 14.960 108.110 15.210 ;
        RECT 107.860 11.350 108.110 11.600 ;
        RECT 107.860 7.740 108.110 7.990 ;
        RECT 107.860 4.130 108.110 4.380 ;
        RECT 107.860 0.520 108.110 0.770 ;
        RECT 107.860 -3.090 108.110 -2.840 ;
        RECT 107.860 -6.700 108.110 -6.450 ;
        RECT 107.860 -10.310 108.110 -10.060 ;
        RECT 107.860 -13.920 108.110 -13.670 ;
        RECT 107.860 -17.530 108.110 -17.280 ;
        RECT 107.860 -21.140 108.110 -20.890 ;
        RECT 107.860 -24.750 108.110 -24.500 ;
        RECT 107.860 -28.360 108.110 -28.110 ;
        RECT 107.860 -31.970 108.110 -31.720 ;
        RECT 107.860 -35.580 108.110 -35.330 ;
        RECT 107.860 -39.190 108.110 -38.940 ;
      LAYER met1 ;
        RECT 107.650 -43.100 108.330 19.120 ;
    END
  END BLb15
  PIN WL0
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER li1 ;
        RECT 7.340 16.220 7.790 16.670 ;
        RECT 20.840 16.220 21.290 16.670 ;
        RECT 34.340 16.220 34.790 16.670 ;
        RECT 47.840 16.220 48.290 16.670 ;
        RECT 61.340 16.220 61.790 16.670 ;
        RECT 74.840 16.220 75.290 16.670 ;
        RECT 88.340 16.220 88.790 16.670 ;
        RECT 101.840 16.220 102.290 16.670 ;
        RECT 115.340 16.220 115.790 16.670 ;
        RECT 128.840 16.220 129.290 16.670 ;
        RECT 142.340 16.220 142.790 16.670 ;
        RECT 155.840 16.220 156.290 16.670 ;
        RECT 169.340 16.220 169.790 16.670 ;
        RECT 182.840 16.220 183.290 16.670 ;
        RECT 196.340 16.220 196.790 16.670 ;
        RECT 209.840 16.220 210.290 16.670 ;
        RECT 0.590 15.310 1.040 15.750 ;
        RECT 14.090 15.310 14.540 15.750 ;
        RECT 27.590 15.310 28.040 15.750 ;
        RECT 41.090 15.310 41.540 15.750 ;
        RECT 54.590 15.310 55.040 15.750 ;
        RECT 68.090 15.310 68.540 15.750 ;
        RECT 81.590 15.310 82.040 15.750 ;
        RECT 95.090 15.310 95.540 15.750 ;
        RECT 108.590 15.310 109.040 15.750 ;
        RECT 122.090 15.310 122.540 15.750 ;
        RECT 135.590 15.310 136.040 15.750 ;
        RECT 149.090 15.310 149.540 15.750 ;
        RECT 162.590 15.310 163.040 15.750 ;
        RECT 176.090 15.310 176.540 15.750 ;
        RECT 189.590 15.310 190.040 15.750 ;
        RECT 203.090 15.310 203.540 15.750 ;
        RECT 216.590 15.310 217.040 15.750 ;
      LAYER mcon ;
        RECT 7.440 16.320 7.690 16.570 ;
        RECT 20.940 16.320 21.190 16.570 ;
        RECT 34.440 16.320 34.690 16.570 ;
        RECT 47.940 16.320 48.190 16.570 ;
        RECT 61.440 16.320 61.690 16.570 ;
        RECT 74.940 16.320 75.190 16.570 ;
        RECT 88.440 16.320 88.690 16.570 ;
        RECT 101.940 16.320 102.190 16.570 ;
        RECT 115.440 16.320 115.690 16.570 ;
        RECT 128.940 16.320 129.190 16.570 ;
        RECT 142.440 16.320 142.690 16.570 ;
        RECT 155.940 16.320 156.190 16.570 ;
        RECT 169.440 16.320 169.690 16.570 ;
        RECT 182.940 16.320 183.190 16.570 ;
        RECT 196.440 16.320 196.690 16.570 ;
        RECT 209.940 16.320 210.190 16.570 ;
        RECT 0.680 15.400 0.950 15.670 ;
        RECT 14.180 15.400 14.450 15.670 ;
        RECT 27.680 15.400 27.950 15.670 ;
        RECT 41.180 15.400 41.450 15.670 ;
        RECT 54.680 15.400 54.950 15.670 ;
        RECT 68.180 15.400 68.450 15.670 ;
        RECT 81.680 15.400 81.950 15.670 ;
        RECT 95.180 15.400 95.450 15.670 ;
        RECT 108.680 15.400 108.950 15.670 ;
        RECT 122.180 15.400 122.450 15.670 ;
        RECT 135.680 15.400 135.950 15.670 ;
        RECT 149.180 15.400 149.450 15.670 ;
        RECT 162.680 15.400 162.950 15.670 ;
        RECT 176.180 15.400 176.450 15.670 ;
        RECT 189.680 15.400 189.950 15.670 ;
        RECT 203.180 15.400 203.450 15.670 ;
        RECT 216.680 15.400 216.950 15.670 ;
      LAYER met1 ;
        RECT 0.590 15.760 1.050 16.230 ;
        RECT 0.580 15.750 1.050 15.760 ;
        RECT 7.330 15.750 7.800 16.680 ;
        RECT 0.580 15.310 1.040 15.750 ;
        RECT 14.080 15.310 14.550 16.230 ;
        RECT 20.830 15.750 21.300 16.680 ;
        RECT 27.580 15.310 28.050 16.230 ;
        RECT 34.330 15.750 34.800 16.680 ;
        RECT 41.080 15.310 41.550 16.230 ;
        RECT 47.830 15.750 48.300 16.680 ;
        RECT 54.580 15.310 55.050 16.230 ;
        RECT 61.330 15.750 61.800 16.680 ;
        RECT 68.080 15.310 68.550 16.230 ;
        RECT 74.830 15.750 75.300 16.680 ;
        RECT 81.580 15.310 82.050 16.230 ;
        RECT 88.330 15.750 88.800 16.680 ;
        RECT 95.080 15.310 95.550 16.230 ;
        RECT 101.830 15.750 102.300 16.680 ;
        RECT 108.580 15.310 109.050 16.230 ;
        RECT 115.330 15.750 115.800 16.680 ;
        RECT 122.080 15.310 122.550 16.230 ;
        RECT 128.830 15.750 129.300 16.680 ;
        RECT 135.580 15.310 136.050 16.230 ;
        RECT 142.330 15.750 142.800 16.680 ;
        RECT 149.080 15.310 149.550 16.230 ;
        RECT 155.830 15.750 156.300 16.680 ;
        RECT 162.580 15.310 163.050 16.230 ;
        RECT 169.330 15.750 169.800 16.680 ;
        RECT 176.080 15.310 176.550 16.230 ;
        RECT 182.830 15.750 183.300 16.680 ;
        RECT 189.580 15.310 190.050 16.230 ;
        RECT 196.330 15.750 196.800 16.680 ;
        RECT 203.080 15.310 203.550 16.230 ;
        RECT 209.830 15.750 210.300 16.680 ;
        RECT 216.580 15.760 217.040 16.230 ;
        RECT 216.580 15.750 217.050 15.760 ;
        RECT 216.590 15.310 217.050 15.750 ;
      LAYER via ;
        RECT 0.680 15.900 0.950 16.170 ;
        RECT 7.430 15.880 7.700 16.150 ;
        RECT 14.180 15.900 14.450 16.170 ;
        RECT 20.930 15.880 21.200 16.150 ;
        RECT 27.680 15.900 27.950 16.170 ;
        RECT 34.430 15.880 34.700 16.150 ;
        RECT 41.180 15.900 41.450 16.170 ;
        RECT 47.930 15.880 48.200 16.150 ;
        RECT 54.680 15.900 54.950 16.170 ;
        RECT 61.430 15.880 61.700 16.150 ;
        RECT 68.180 15.900 68.450 16.170 ;
        RECT 74.930 15.880 75.200 16.150 ;
        RECT 81.680 15.900 81.950 16.170 ;
        RECT 88.430 15.880 88.700 16.150 ;
        RECT 95.180 15.900 95.450 16.170 ;
        RECT 101.930 15.880 102.200 16.150 ;
        RECT 108.680 15.900 108.950 16.170 ;
        RECT 115.430 15.880 115.700 16.150 ;
        RECT 122.180 15.900 122.450 16.170 ;
        RECT 128.930 15.880 129.200 16.150 ;
        RECT 135.680 15.900 135.950 16.170 ;
        RECT 142.430 15.880 142.700 16.150 ;
        RECT 149.180 15.900 149.450 16.170 ;
        RECT 155.930 15.880 156.200 16.150 ;
        RECT 162.680 15.900 162.950 16.170 ;
        RECT 169.430 15.880 169.700 16.150 ;
        RECT 176.180 15.900 176.450 16.170 ;
        RECT 182.930 15.880 183.200 16.150 ;
        RECT 189.680 15.900 189.950 16.170 ;
        RECT 196.430 15.880 196.700 16.150 ;
        RECT 203.180 15.900 203.450 16.170 ;
        RECT 209.930 15.880 210.200 16.150 ;
        RECT 216.680 15.900 216.950 16.170 ;
      LAYER met2 ;
        RECT 0.580 15.760 217.050 16.270 ;
        RECT 0.590 15.750 217.040 15.760 ;
    END
  END WL0
  PIN WL1
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER li1 ;
        RECT 0.590 14.420 1.040 14.860 ;
        RECT 14.090 14.420 14.540 14.860 ;
        RECT 27.590 14.420 28.040 14.860 ;
        RECT 41.090 14.420 41.540 14.860 ;
        RECT 54.590 14.420 55.040 14.860 ;
        RECT 68.090 14.420 68.540 14.860 ;
        RECT 81.590 14.420 82.040 14.860 ;
        RECT 95.090 14.420 95.540 14.860 ;
        RECT 108.590 14.420 109.040 14.860 ;
        RECT 122.090 14.420 122.540 14.860 ;
        RECT 135.590 14.420 136.040 14.860 ;
        RECT 149.090 14.420 149.540 14.860 ;
        RECT 162.590 14.420 163.040 14.860 ;
        RECT 176.090 14.420 176.540 14.860 ;
        RECT 189.590 14.420 190.040 14.860 ;
        RECT 203.090 14.420 203.540 14.860 ;
        RECT 216.590 14.420 217.040 14.860 ;
        RECT 7.340 13.500 7.790 13.950 ;
        RECT 20.840 13.500 21.290 13.950 ;
        RECT 34.340 13.500 34.790 13.950 ;
        RECT 47.840 13.500 48.290 13.950 ;
        RECT 61.340 13.500 61.790 13.950 ;
        RECT 74.840 13.500 75.290 13.950 ;
        RECT 88.340 13.500 88.790 13.950 ;
        RECT 101.840 13.500 102.290 13.950 ;
        RECT 115.340 13.500 115.790 13.950 ;
        RECT 128.840 13.500 129.290 13.950 ;
        RECT 142.340 13.500 142.790 13.950 ;
        RECT 155.840 13.500 156.290 13.950 ;
        RECT 169.340 13.500 169.790 13.950 ;
        RECT 182.840 13.500 183.290 13.950 ;
        RECT 196.340 13.500 196.790 13.950 ;
        RECT 209.840 13.500 210.290 13.950 ;
      LAYER mcon ;
        RECT 0.680 14.500 0.950 14.770 ;
        RECT 14.180 14.500 14.450 14.770 ;
        RECT 27.680 14.500 27.950 14.770 ;
        RECT 41.180 14.500 41.450 14.770 ;
        RECT 54.680 14.500 54.950 14.770 ;
        RECT 68.180 14.500 68.450 14.770 ;
        RECT 81.680 14.500 81.950 14.770 ;
        RECT 95.180 14.500 95.450 14.770 ;
        RECT 108.680 14.500 108.950 14.770 ;
        RECT 122.180 14.500 122.450 14.770 ;
        RECT 135.680 14.500 135.950 14.770 ;
        RECT 149.180 14.500 149.450 14.770 ;
        RECT 162.680 14.500 162.950 14.770 ;
        RECT 176.180 14.500 176.450 14.770 ;
        RECT 189.680 14.500 189.950 14.770 ;
        RECT 203.180 14.500 203.450 14.770 ;
        RECT 216.680 14.500 216.950 14.770 ;
        RECT 7.440 13.600 7.690 13.850 ;
        RECT 20.940 13.600 21.190 13.850 ;
        RECT 34.440 13.600 34.690 13.850 ;
        RECT 47.940 13.600 48.190 13.850 ;
        RECT 61.440 13.600 61.690 13.850 ;
        RECT 74.940 13.600 75.190 13.850 ;
        RECT 88.440 13.600 88.690 13.850 ;
        RECT 101.940 13.600 102.190 13.850 ;
        RECT 115.440 13.600 115.690 13.850 ;
        RECT 128.940 13.600 129.190 13.850 ;
        RECT 142.440 13.600 142.690 13.850 ;
        RECT 155.940 13.600 156.190 13.850 ;
        RECT 169.440 13.600 169.690 13.850 ;
        RECT 182.940 13.600 183.190 13.850 ;
        RECT 196.440 13.600 196.690 13.850 ;
        RECT 209.940 13.600 210.190 13.850 ;
      LAYER met1 ;
        RECT 0.580 14.420 1.040 14.860 ;
        RECT 0.580 14.410 1.050 14.420 ;
        RECT 0.590 13.940 1.050 14.410 ;
        RECT 7.330 13.490 7.800 14.420 ;
        RECT 14.080 13.940 14.550 14.860 ;
        RECT 20.830 13.490 21.300 14.420 ;
        RECT 27.580 13.940 28.050 14.860 ;
        RECT 34.330 13.490 34.800 14.420 ;
        RECT 41.080 13.940 41.550 14.860 ;
        RECT 47.830 13.490 48.300 14.420 ;
        RECT 54.580 13.940 55.050 14.860 ;
        RECT 61.330 13.490 61.800 14.420 ;
        RECT 68.080 13.940 68.550 14.860 ;
        RECT 74.830 13.490 75.300 14.420 ;
        RECT 81.580 13.940 82.050 14.860 ;
        RECT 88.330 13.490 88.800 14.420 ;
        RECT 95.080 13.940 95.550 14.860 ;
        RECT 101.830 13.490 102.300 14.420 ;
        RECT 108.580 13.940 109.050 14.860 ;
        RECT 115.330 13.490 115.800 14.420 ;
        RECT 122.080 13.940 122.550 14.860 ;
        RECT 128.830 13.490 129.300 14.420 ;
        RECT 135.580 13.940 136.050 14.860 ;
        RECT 142.330 13.490 142.800 14.420 ;
        RECT 149.080 13.940 149.550 14.860 ;
        RECT 155.830 13.490 156.300 14.420 ;
        RECT 162.580 13.940 163.050 14.860 ;
        RECT 169.330 13.490 169.800 14.420 ;
        RECT 176.080 13.940 176.550 14.860 ;
        RECT 182.830 13.490 183.300 14.420 ;
        RECT 189.580 13.940 190.050 14.860 ;
        RECT 196.330 13.490 196.800 14.420 ;
        RECT 203.080 13.940 203.550 14.860 ;
        RECT 216.590 14.420 217.050 14.860 ;
        RECT 209.830 13.490 210.300 14.420 ;
        RECT 216.580 14.410 217.050 14.420 ;
        RECT 216.580 13.940 217.040 14.410 ;
      LAYER via ;
        RECT 0.680 14.000 0.950 14.270 ;
        RECT 7.430 14.050 7.700 14.320 ;
        RECT 14.180 14.000 14.450 14.270 ;
        RECT 20.930 14.050 21.200 14.320 ;
        RECT 27.680 14.000 27.950 14.270 ;
        RECT 34.430 14.050 34.700 14.320 ;
        RECT 41.180 14.000 41.450 14.270 ;
        RECT 47.930 14.050 48.200 14.320 ;
        RECT 54.680 14.000 54.950 14.270 ;
        RECT 61.430 14.050 61.700 14.320 ;
        RECT 68.180 14.000 68.450 14.270 ;
        RECT 74.930 14.050 75.200 14.320 ;
        RECT 81.680 14.000 81.950 14.270 ;
        RECT 88.430 14.050 88.700 14.320 ;
        RECT 95.180 14.000 95.450 14.270 ;
        RECT 101.930 14.050 102.200 14.320 ;
        RECT 108.680 14.000 108.950 14.270 ;
        RECT 115.430 14.050 115.700 14.320 ;
        RECT 122.180 14.000 122.450 14.270 ;
        RECT 128.930 14.050 129.200 14.320 ;
        RECT 135.680 14.000 135.950 14.270 ;
        RECT 142.430 14.050 142.700 14.320 ;
        RECT 149.180 14.000 149.450 14.270 ;
        RECT 155.930 14.050 156.200 14.320 ;
        RECT 162.680 14.000 162.950 14.270 ;
        RECT 169.430 14.050 169.700 14.320 ;
        RECT 176.180 14.000 176.450 14.270 ;
        RECT 182.930 14.050 183.200 14.320 ;
        RECT 189.680 14.000 189.950 14.270 ;
        RECT 196.430 14.050 196.700 14.320 ;
        RECT 203.180 14.000 203.450 14.270 ;
        RECT 209.930 14.050 210.200 14.320 ;
        RECT 216.680 14.000 216.950 14.270 ;
      LAYER met2 ;
        RECT 0.590 13.910 217.040 14.430 ;
        RECT 0.590 13.900 1.070 13.910 ;
        RECT 108.560 13.900 109.070 13.910 ;
        RECT 216.560 13.900 217.040 13.910 ;
    END
  END WL1
  PIN WL2
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER li1 ;
        RECT 7.340 12.610 7.790 13.060 ;
        RECT 20.840 12.610 21.290 13.060 ;
        RECT 34.340 12.610 34.790 13.060 ;
        RECT 47.840 12.610 48.290 13.060 ;
        RECT 61.340 12.610 61.790 13.060 ;
        RECT 74.840 12.610 75.290 13.060 ;
        RECT 88.340 12.610 88.790 13.060 ;
        RECT 101.840 12.610 102.290 13.060 ;
        RECT 115.340 12.610 115.790 13.060 ;
        RECT 128.840 12.610 129.290 13.060 ;
        RECT 142.340 12.610 142.790 13.060 ;
        RECT 155.840 12.610 156.290 13.060 ;
        RECT 169.340 12.610 169.790 13.060 ;
        RECT 182.840 12.610 183.290 13.060 ;
        RECT 196.340 12.610 196.790 13.060 ;
        RECT 209.840 12.610 210.290 13.060 ;
        RECT 0.590 11.700 1.040 12.140 ;
        RECT 14.090 11.700 14.540 12.140 ;
        RECT 27.590 11.700 28.040 12.140 ;
        RECT 41.090 11.700 41.540 12.140 ;
        RECT 54.590 11.700 55.040 12.140 ;
        RECT 68.090 11.700 68.540 12.140 ;
        RECT 81.590 11.700 82.040 12.140 ;
        RECT 95.090 11.700 95.540 12.140 ;
        RECT 108.590 11.700 109.040 12.140 ;
        RECT 122.090 11.700 122.540 12.140 ;
        RECT 135.590 11.700 136.040 12.140 ;
        RECT 149.090 11.700 149.540 12.140 ;
        RECT 162.590 11.700 163.040 12.140 ;
        RECT 176.090 11.700 176.540 12.140 ;
        RECT 189.590 11.700 190.040 12.140 ;
        RECT 203.090 11.700 203.540 12.140 ;
        RECT 216.590 11.700 217.040 12.140 ;
      LAYER mcon ;
        RECT 7.440 12.710 7.690 12.960 ;
        RECT 20.940 12.710 21.190 12.960 ;
        RECT 34.440 12.710 34.690 12.960 ;
        RECT 47.940 12.710 48.190 12.960 ;
        RECT 61.440 12.710 61.690 12.960 ;
        RECT 74.940 12.710 75.190 12.960 ;
        RECT 88.440 12.710 88.690 12.960 ;
        RECT 101.940 12.710 102.190 12.960 ;
        RECT 115.440 12.710 115.690 12.960 ;
        RECT 128.940 12.710 129.190 12.960 ;
        RECT 142.440 12.710 142.690 12.960 ;
        RECT 155.940 12.710 156.190 12.960 ;
        RECT 169.440 12.710 169.690 12.960 ;
        RECT 182.940 12.710 183.190 12.960 ;
        RECT 196.440 12.710 196.690 12.960 ;
        RECT 209.940 12.710 210.190 12.960 ;
        RECT 0.680 11.790 0.950 12.060 ;
        RECT 14.180 11.790 14.450 12.060 ;
        RECT 27.680 11.790 27.950 12.060 ;
        RECT 41.180 11.790 41.450 12.060 ;
        RECT 54.680 11.790 54.950 12.060 ;
        RECT 68.180 11.790 68.450 12.060 ;
        RECT 81.680 11.790 81.950 12.060 ;
        RECT 95.180 11.790 95.450 12.060 ;
        RECT 108.680 11.790 108.950 12.060 ;
        RECT 122.180 11.790 122.450 12.060 ;
        RECT 135.680 11.790 135.950 12.060 ;
        RECT 149.180 11.790 149.450 12.060 ;
        RECT 162.680 11.790 162.950 12.060 ;
        RECT 176.180 11.790 176.450 12.060 ;
        RECT 189.680 11.790 189.950 12.060 ;
        RECT 203.180 11.790 203.450 12.060 ;
        RECT 216.680 11.790 216.950 12.060 ;
      LAYER met1 ;
        RECT 0.590 12.150 1.050 12.620 ;
        RECT 0.580 12.140 1.050 12.150 ;
        RECT 7.330 12.140 7.800 13.070 ;
        RECT 0.580 11.700 1.040 12.140 ;
        RECT 14.080 11.700 14.550 12.620 ;
        RECT 20.830 12.140 21.300 13.070 ;
        RECT 27.580 11.700 28.050 12.620 ;
        RECT 34.330 12.140 34.800 13.070 ;
        RECT 41.080 11.700 41.550 12.620 ;
        RECT 47.830 12.140 48.300 13.070 ;
        RECT 54.580 11.700 55.050 12.620 ;
        RECT 61.330 12.140 61.800 13.070 ;
        RECT 68.080 11.700 68.550 12.620 ;
        RECT 74.830 12.140 75.300 13.070 ;
        RECT 81.580 11.700 82.050 12.620 ;
        RECT 88.330 12.140 88.800 13.070 ;
        RECT 95.080 11.700 95.550 12.620 ;
        RECT 101.830 12.140 102.300 13.070 ;
        RECT 108.580 11.700 109.050 12.620 ;
        RECT 115.330 12.140 115.800 13.070 ;
        RECT 122.080 11.700 122.550 12.620 ;
        RECT 128.830 12.140 129.300 13.070 ;
        RECT 135.580 11.700 136.050 12.620 ;
        RECT 142.330 12.140 142.800 13.070 ;
        RECT 149.080 11.700 149.550 12.620 ;
        RECT 155.830 12.140 156.300 13.070 ;
        RECT 162.580 11.700 163.050 12.620 ;
        RECT 169.330 12.140 169.800 13.070 ;
        RECT 176.080 11.700 176.550 12.620 ;
        RECT 182.830 12.140 183.300 13.070 ;
        RECT 189.580 11.700 190.050 12.620 ;
        RECT 196.330 12.140 196.800 13.070 ;
        RECT 203.080 11.700 203.550 12.620 ;
        RECT 209.830 12.140 210.300 13.070 ;
        RECT 216.580 12.150 217.040 12.620 ;
        RECT 216.580 12.140 217.050 12.150 ;
        RECT 216.590 11.700 217.050 12.140 ;
      LAYER via ;
        RECT 0.680 12.290 0.950 12.560 ;
        RECT 7.430 12.270 7.700 12.540 ;
        RECT 14.180 12.290 14.450 12.560 ;
        RECT 20.930 12.240 21.200 12.510 ;
        RECT 27.680 12.290 27.950 12.560 ;
        RECT 34.430 12.240 34.700 12.510 ;
        RECT 41.180 12.290 41.450 12.560 ;
        RECT 47.930 12.270 48.200 12.540 ;
        RECT 54.680 12.290 54.950 12.560 ;
        RECT 61.430 12.270 61.700 12.540 ;
        RECT 68.180 12.290 68.450 12.560 ;
        RECT 74.930 12.240 75.200 12.510 ;
        RECT 81.680 12.290 81.950 12.560 ;
        RECT 88.430 12.240 88.700 12.510 ;
        RECT 95.180 12.290 95.450 12.560 ;
        RECT 101.930 12.270 102.200 12.540 ;
        RECT 108.680 12.290 108.950 12.560 ;
        RECT 115.430 12.270 115.700 12.540 ;
        RECT 122.180 12.290 122.450 12.560 ;
        RECT 128.930 12.240 129.200 12.510 ;
        RECT 135.680 12.290 135.950 12.560 ;
        RECT 142.430 12.240 142.700 12.510 ;
        RECT 149.180 12.290 149.450 12.560 ;
        RECT 155.930 12.270 156.200 12.540 ;
        RECT 162.680 12.290 162.950 12.560 ;
        RECT 169.430 12.270 169.700 12.540 ;
        RECT 176.180 12.290 176.450 12.560 ;
        RECT 182.930 12.240 183.200 12.510 ;
        RECT 189.680 12.290 189.950 12.560 ;
        RECT 196.430 12.240 196.700 12.510 ;
        RECT 203.180 12.290 203.450 12.560 ;
        RECT 209.930 12.270 210.200 12.540 ;
        RECT 216.680 12.290 216.950 12.560 ;
      LAYER met2 ;
        RECT 0.590 12.660 1.070 12.670 ;
        RECT 108.560 12.660 109.070 12.670 ;
        RECT 216.560 12.660 217.040 12.670 ;
        RECT 0.590 12.650 14.590 12.660 ;
        RECT 41.040 12.650 68.590 12.660 ;
        RECT 95.040 12.650 122.590 12.660 ;
        RECT 149.040 12.650 176.590 12.660 ;
        RECT 203.040 12.650 217.040 12.660 ;
        RECT 0.590 12.630 217.040 12.650 ;
        RECT 0.580 12.150 217.050 12.630 ;
        RECT 0.590 12.140 217.040 12.150 ;
        RECT 14.040 12.130 41.590 12.140 ;
        RECT 68.040 12.130 95.590 12.140 ;
        RECT 122.040 12.130 149.590 12.140 ;
        RECT 176.040 12.130 203.590 12.140 ;
    END
  END WL2
  PIN WL3
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER li1 ;
        RECT 0.590 10.810 1.040 11.250 ;
        RECT 14.090 10.810 14.540 11.250 ;
        RECT 27.590 10.810 28.040 11.250 ;
        RECT 41.090 10.810 41.540 11.250 ;
        RECT 54.590 10.810 55.040 11.250 ;
        RECT 68.090 10.810 68.540 11.250 ;
        RECT 81.590 10.810 82.040 11.250 ;
        RECT 95.090 10.810 95.540 11.250 ;
        RECT 108.590 10.810 109.040 11.250 ;
        RECT 122.090 10.810 122.540 11.250 ;
        RECT 135.590 10.810 136.040 11.250 ;
        RECT 149.090 10.810 149.540 11.250 ;
        RECT 162.590 10.810 163.040 11.250 ;
        RECT 176.090 10.810 176.540 11.250 ;
        RECT 189.590 10.810 190.040 11.250 ;
        RECT 203.090 10.810 203.540 11.250 ;
        RECT 216.590 10.810 217.040 11.250 ;
        RECT 7.340 9.890 7.790 10.340 ;
        RECT 20.840 9.890 21.290 10.340 ;
        RECT 34.340 9.890 34.790 10.340 ;
        RECT 47.840 9.890 48.290 10.340 ;
        RECT 61.340 9.890 61.790 10.340 ;
        RECT 74.840 9.890 75.290 10.340 ;
        RECT 88.340 9.890 88.790 10.340 ;
        RECT 101.840 9.890 102.290 10.340 ;
        RECT 115.340 9.890 115.790 10.340 ;
        RECT 128.840 9.890 129.290 10.340 ;
        RECT 142.340 9.890 142.790 10.340 ;
        RECT 155.840 9.890 156.290 10.340 ;
        RECT 169.340 9.890 169.790 10.340 ;
        RECT 182.840 9.890 183.290 10.340 ;
        RECT 196.340 9.890 196.790 10.340 ;
        RECT 209.840 9.890 210.290 10.340 ;
      LAYER mcon ;
        RECT 0.680 10.890 0.950 11.160 ;
        RECT 14.180 10.890 14.450 11.160 ;
        RECT 27.680 10.890 27.950 11.160 ;
        RECT 41.180 10.890 41.450 11.160 ;
        RECT 54.680 10.890 54.950 11.160 ;
        RECT 68.180 10.890 68.450 11.160 ;
        RECT 81.680 10.890 81.950 11.160 ;
        RECT 95.180 10.890 95.450 11.160 ;
        RECT 108.680 10.890 108.950 11.160 ;
        RECT 122.180 10.890 122.450 11.160 ;
        RECT 135.680 10.890 135.950 11.160 ;
        RECT 149.180 10.890 149.450 11.160 ;
        RECT 162.680 10.890 162.950 11.160 ;
        RECT 176.180 10.890 176.450 11.160 ;
        RECT 189.680 10.890 189.950 11.160 ;
        RECT 203.180 10.890 203.450 11.160 ;
        RECT 216.680 10.890 216.950 11.160 ;
        RECT 7.440 9.990 7.690 10.240 ;
        RECT 20.940 9.990 21.190 10.240 ;
        RECT 34.440 9.990 34.690 10.240 ;
        RECT 47.940 9.990 48.190 10.240 ;
        RECT 61.440 9.990 61.690 10.240 ;
        RECT 74.940 9.990 75.190 10.240 ;
        RECT 88.440 9.990 88.690 10.240 ;
        RECT 101.940 9.990 102.190 10.240 ;
        RECT 115.440 9.990 115.690 10.240 ;
        RECT 128.940 9.990 129.190 10.240 ;
        RECT 142.440 9.990 142.690 10.240 ;
        RECT 155.940 9.990 156.190 10.240 ;
        RECT 169.440 9.990 169.690 10.240 ;
        RECT 182.940 9.990 183.190 10.240 ;
        RECT 196.440 9.990 196.690 10.240 ;
        RECT 209.940 9.990 210.190 10.240 ;
      LAYER met1 ;
        RECT 0.580 10.810 1.040 11.250 ;
        RECT 0.580 10.800 1.050 10.810 ;
        RECT 0.590 10.330 1.050 10.800 ;
        RECT 7.330 9.880 7.800 10.810 ;
        RECT 14.080 10.330 14.550 11.250 ;
        RECT 20.830 9.880 21.300 10.810 ;
        RECT 27.580 10.330 28.050 11.250 ;
        RECT 34.330 9.880 34.800 10.810 ;
        RECT 41.080 10.330 41.550 11.250 ;
        RECT 47.830 9.880 48.300 10.810 ;
        RECT 54.580 10.330 55.050 11.250 ;
        RECT 61.330 9.880 61.800 10.810 ;
        RECT 68.080 10.330 68.550 11.250 ;
        RECT 74.830 9.880 75.300 10.810 ;
        RECT 81.580 10.330 82.050 11.250 ;
        RECT 88.330 9.880 88.800 10.810 ;
        RECT 95.080 10.330 95.550 11.250 ;
        RECT 101.830 9.880 102.300 10.810 ;
        RECT 108.580 10.330 109.050 11.250 ;
        RECT 115.330 9.880 115.800 10.810 ;
        RECT 122.080 10.330 122.550 11.250 ;
        RECT 128.830 9.880 129.300 10.810 ;
        RECT 135.580 10.330 136.050 11.250 ;
        RECT 142.330 9.880 142.800 10.810 ;
        RECT 149.080 10.330 149.550 11.250 ;
        RECT 155.830 9.880 156.300 10.810 ;
        RECT 162.580 10.330 163.050 11.250 ;
        RECT 169.330 9.880 169.800 10.810 ;
        RECT 176.080 10.330 176.550 11.250 ;
        RECT 182.830 9.880 183.300 10.810 ;
        RECT 189.580 10.330 190.050 11.250 ;
        RECT 196.330 9.880 196.800 10.810 ;
        RECT 203.080 10.330 203.550 11.250 ;
        RECT 216.590 10.810 217.050 11.250 ;
        RECT 209.830 9.880 210.300 10.810 ;
        RECT 216.580 10.800 217.050 10.810 ;
        RECT 216.580 10.330 217.040 10.800 ;
      LAYER via ;
        RECT 0.680 10.390 0.950 10.660 ;
        RECT 7.430 10.440 7.700 10.710 ;
        RECT 14.180 10.390 14.450 10.660 ;
        RECT 20.930 10.410 21.200 10.680 ;
        RECT 27.680 10.390 27.950 10.660 ;
        RECT 34.430 10.410 34.700 10.680 ;
        RECT 41.180 10.390 41.450 10.660 ;
        RECT 47.930 10.440 48.200 10.710 ;
        RECT 54.680 10.390 54.950 10.660 ;
        RECT 61.430 10.440 61.700 10.710 ;
        RECT 68.180 10.390 68.450 10.660 ;
        RECT 74.930 10.410 75.200 10.680 ;
        RECT 81.680 10.390 81.950 10.660 ;
        RECT 88.430 10.410 88.700 10.680 ;
        RECT 95.180 10.390 95.450 10.660 ;
        RECT 101.930 10.440 102.200 10.710 ;
        RECT 108.680 10.390 108.950 10.660 ;
        RECT 115.430 10.440 115.700 10.710 ;
        RECT 122.180 10.390 122.450 10.660 ;
        RECT 128.930 10.410 129.200 10.680 ;
        RECT 135.680 10.390 135.950 10.660 ;
        RECT 142.430 10.410 142.700 10.680 ;
        RECT 149.180 10.390 149.450 10.660 ;
        RECT 155.930 10.440 156.200 10.710 ;
        RECT 162.680 10.390 162.950 10.660 ;
        RECT 169.430 10.440 169.700 10.710 ;
        RECT 176.180 10.390 176.450 10.660 ;
        RECT 182.930 10.410 183.200 10.680 ;
        RECT 189.680 10.390 189.950 10.660 ;
        RECT 196.430 10.410 196.700 10.680 ;
        RECT 203.180 10.390 203.450 10.660 ;
        RECT 209.930 10.440 210.200 10.710 ;
        RECT 216.680 10.390 216.950 10.660 ;
      LAYER met2 ;
        RECT 0.590 10.810 14.590 10.820 ;
        RECT 41.040 10.810 68.590 10.820 ;
        RECT 95.040 10.810 122.590 10.820 ;
        RECT 149.040 10.810 176.590 10.820 ;
        RECT 203.040 10.810 217.040 10.820 ;
        RECT 0.590 10.790 217.040 10.810 ;
        RECT 0.580 10.310 217.050 10.790 ;
        RECT 0.590 10.300 217.040 10.310 ;
        RECT 14.040 10.290 41.590 10.300 ;
        RECT 68.040 10.290 95.590 10.300 ;
        RECT 122.040 10.290 149.590 10.300 ;
        RECT 176.040 10.290 203.590 10.300 ;
    END
  END WL3
  PIN WL4
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER li1 ;
        RECT 7.340 9.000 7.790 9.450 ;
        RECT 20.840 9.000 21.290 9.450 ;
        RECT 34.340 9.000 34.790 9.450 ;
        RECT 47.840 9.000 48.290 9.450 ;
        RECT 61.340 9.000 61.790 9.450 ;
        RECT 74.840 9.000 75.290 9.450 ;
        RECT 88.340 9.000 88.790 9.450 ;
        RECT 101.840 9.000 102.290 9.450 ;
        RECT 115.340 9.000 115.790 9.450 ;
        RECT 128.840 9.000 129.290 9.450 ;
        RECT 142.340 9.000 142.790 9.450 ;
        RECT 155.840 9.000 156.290 9.450 ;
        RECT 169.340 9.000 169.790 9.450 ;
        RECT 182.840 9.000 183.290 9.450 ;
        RECT 196.340 9.000 196.790 9.450 ;
        RECT 209.840 9.000 210.290 9.450 ;
        RECT 0.590 8.090 1.040 8.530 ;
        RECT 14.090 8.090 14.540 8.530 ;
        RECT 27.590 8.090 28.040 8.530 ;
        RECT 41.090 8.090 41.540 8.530 ;
        RECT 54.590 8.090 55.040 8.530 ;
        RECT 68.090 8.090 68.540 8.530 ;
        RECT 81.590 8.090 82.040 8.530 ;
        RECT 95.090 8.090 95.540 8.530 ;
        RECT 108.590 8.090 109.040 8.530 ;
        RECT 122.090 8.090 122.540 8.530 ;
        RECT 135.590 8.090 136.040 8.530 ;
        RECT 149.090 8.090 149.540 8.530 ;
        RECT 162.590 8.090 163.040 8.530 ;
        RECT 176.090 8.090 176.540 8.530 ;
        RECT 189.590 8.090 190.040 8.530 ;
        RECT 203.090 8.090 203.540 8.530 ;
        RECT 216.590 8.090 217.040 8.530 ;
      LAYER mcon ;
        RECT 7.440 9.100 7.690 9.350 ;
        RECT 20.940 9.100 21.190 9.350 ;
        RECT 34.440 9.100 34.690 9.350 ;
        RECT 47.940 9.100 48.190 9.350 ;
        RECT 61.440 9.100 61.690 9.350 ;
        RECT 74.940 9.100 75.190 9.350 ;
        RECT 88.440 9.100 88.690 9.350 ;
        RECT 101.940 9.100 102.190 9.350 ;
        RECT 115.440 9.100 115.690 9.350 ;
        RECT 128.940 9.100 129.190 9.350 ;
        RECT 142.440 9.100 142.690 9.350 ;
        RECT 155.940 9.100 156.190 9.350 ;
        RECT 169.440 9.100 169.690 9.350 ;
        RECT 182.940 9.100 183.190 9.350 ;
        RECT 196.440 9.100 196.690 9.350 ;
        RECT 209.940 9.100 210.190 9.350 ;
        RECT 0.680 8.180 0.950 8.450 ;
        RECT 14.180 8.180 14.450 8.450 ;
        RECT 27.680 8.180 27.950 8.450 ;
        RECT 41.180 8.180 41.450 8.450 ;
        RECT 54.680 8.180 54.950 8.450 ;
        RECT 68.180 8.180 68.450 8.450 ;
        RECT 81.680 8.180 81.950 8.450 ;
        RECT 95.180 8.180 95.450 8.450 ;
        RECT 108.680 8.180 108.950 8.450 ;
        RECT 122.180 8.180 122.450 8.450 ;
        RECT 135.680 8.180 135.950 8.450 ;
        RECT 149.180 8.180 149.450 8.450 ;
        RECT 162.680 8.180 162.950 8.450 ;
        RECT 176.180 8.180 176.450 8.450 ;
        RECT 189.680 8.180 189.950 8.450 ;
        RECT 203.180 8.180 203.450 8.450 ;
        RECT 216.680 8.180 216.950 8.450 ;
      LAYER met1 ;
        RECT 0.590 8.540 1.050 9.010 ;
        RECT 0.580 8.530 1.050 8.540 ;
        RECT 7.330 8.530 7.800 9.460 ;
        RECT 0.580 8.090 1.040 8.530 ;
        RECT 14.080 8.090 14.550 9.010 ;
        RECT 20.830 8.530 21.300 9.460 ;
        RECT 27.580 8.090 28.050 9.010 ;
        RECT 34.330 8.530 34.800 9.460 ;
        RECT 41.080 8.090 41.550 9.010 ;
        RECT 47.830 8.530 48.300 9.460 ;
        RECT 54.580 8.090 55.050 9.010 ;
        RECT 61.330 8.530 61.800 9.460 ;
        RECT 68.080 8.090 68.550 9.010 ;
        RECT 74.830 8.530 75.300 9.460 ;
        RECT 81.580 8.090 82.050 9.010 ;
        RECT 88.330 8.530 88.800 9.460 ;
        RECT 95.080 8.090 95.550 9.010 ;
        RECT 101.830 8.530 102.300 9.460 ;
        RECT 108.580 8.090 109.050 9.010 ;
        RECT 115.330 8.530 115.800 9.460 ;
        RECT 122.080 8.090 122.550 9.010 ;
        RECT 128.830 8.530 129.300 9.460 ;
        RECT 135.580 8.090 136.050 9.010 ;
        RECT 142.330 8.530 142.800 9.460 ;
        RECT 149.080 8.090 149.550 9.010 ;
        RECT 155.830 8.530 156.300 9.460 ;
        RECT 162.580 8.090 163.050 9.010 ;
        RECT 169.330 8.530 169.800 9.460 ;
        RECT 176.080 8.090 176.550 9.010 ;
        RECT 182.830 8.530 183.300 9.460 ;
        RECT 189.580 8.090 190.050 9.010 ;
        RECT 196.330 8.530 196.800 9.460 ;
        RECT 203.080 8.090 203.550 9.010 ;
        RECT 209.830 8.530 210.300 9.460 ;
        RECT 216.580 8.540 217.040 9.010 ;
        RECT 216.580 8.530 217.050 8.540 ;
        RECT 216.590 8.090 217.050 8.530 ;
      LAYER via ;
        RECT 0.680 8.680 0.950 8.950 ;
        RECT 7.430 8.630 7.700 8.900 ;
        RECT 14.180 8.680 14.450 8.950 ;
        RECT 20.930 8.660 21.200 8.930 ;
        RECT 27.680 8.680 27.950 8.950 ;
        RECT 34.430 8.660 34.700 8.930 ;
        RECT 41.180 8.680 41.450 8.950 ;
        RECT 47.930 8.630 48.200 8.900 ;
        RECT 54.680 8.680 54.950 8.950 ;
        RECT 61.430 8.630 61.700 8.900 ;
        RECT 68.180 8.680 68.450 8.950 ;
        RECT 74.930 8.660 75.200 8.930 ;
        RECT 81.680 8.680 81.950 8.950 ;
        RECT 88.430 8.660 88.700 8.930 ;
        RECT 95.180 8.680 95.450 8.950 ;
        RECT 101.930 8.630 102.200 8.900 ;
        RECT 108.680 8.680 108.950 8.950 ;
        RECT 115.430 8.630 115.700 8.900 ;
        RECT 122.180 8.680 122.450 8.950 ;
        RECT 128.930 8.660 129.200 8.930 ;
        RECT 135.680 8.680 135.950 8.950 ;
        RECT 142.430 8.660 142.700 8.930 ;
        RECT 149.180 8.680 149.450 8.950 ;
        RECT 155.930 8.630 156.200 8.900 ;
        RECT 162.680 8.680 162.950 8.950 ;
        RECT 169.430 8.630 169.700 8.900 ;
        RECT 176.180 8.680 176.450 8.950 ;
        RECT 182.930 8.660 183.200 8.930 ;
        RECT 189.680 8.680 189.950 8.950 ;
        RECT 196.430 8.660 196.700 8.930 ;
        RECT 203.180 8.680 203.450 8.950 ;
        RECT 209.930 8.630 210.200 8.900 ;
        RECT 216.680 8.680 216.950 8.950 ;
      LAYER met2 ;
        RECT 0.580 9.040 1.060 9.050 ;
        RECT 14.040 9.040 41.590 9.050 ;
        RECT 68.040 9.040 95.590 9.050 ;
        RECT 108.570 9.040 109.060 9.050 ;
        RECT 122.040 9.040 149.590 9.050 ;
        RECT 176.040 9.040 203.590 9.050 ;
        RECT 216.570 9.040 217.050 9.050 ;
        RECT 0.580 8.540 217.050 9.040 ;
        RECT 0.590 8.530 217.040 8.540 ;
        RECT 0.590 8.520 14.590 8.530 ;
        RECT 41.040 8.520 68.590 8.530 ;
        RECT 95.040 8.520 122.590 8.530 ;
        RECT 149.040 8.520 176.590 8.530 ;
        RECT 203.040 8.520 217.040 8.530 ;
    END
  END WL4
  PIN WL5
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER li1 ;
        RECT 0.590 7.200 1.040 7.640 ;
        RECT 14.090 7.200 14.540 7.640 ;
        RECT 27.590 7.200 28.040 7.640 ;
        RECT 41.090 7.200 41.540 7.640 ;
        RECT 54.590 7.200 55.040 7.640 ;
        RECT 68.090 7.200 68.540 7.640 ;
        RECT 81.590 7.200 82.040 7.640 ;
        RECT 95.090 7.200 95.540 7.640 ;
        RECT 108.590 7.200 109.040 7.640 ;
        RECT 122.090 7.200 122.540 7.640 ;
        RECT 135.590 7.200 136.040 7.640 ;
        RECT 149.090 7.200 149.540 7.640 ;
        RECT 162.590 7.200 163.040 7.640 ;
        RECT 176.090 7.200 176.540 7.640 ;
        RECT 189.590 7.200 190.040 7.640 ;
        RECT 203.090 7.200 203.540 7.640 ;
        RECT 216.590 7.200 217.040 7.640 ;
        RECT 7.340 6.280 7.790 6.730 ;
        RECT 20.840 6.280 21.290 6.730 ;
        RECT 34.340 6.280 34.790 6.730 ;
        RECT 47.840 6.280 48.290 6.730 ;
        RECT 61.340 6.280 61.790 6.730 ;
        RECT 74.840 6.280 75.290 6.730 ;
        RECT 88.340 6.280 88.790 6.730 ;
        RECT 101.840 6.280 102.290 6.730 ;
        RECT 115.340 6.280 115.790 6.730 ;
        RECT 128.840 6.280 129.290 6.730 ;
        RECT 142.340 6.280 142.790 6.730 ;
        RECT 155.840 6.280 156.290 6.730 ;
        RECT 169.340 6.280 169.790 6.730 ;
        RECT 182.840 6.280 183.290 6.730 ;
        RECT 196.340 6.280 196.790 6.730 ;
        RECT 209.840 6.280 210.290 6.730 ;
      LAYER mcon ;
        RECT 0.680 7.280 0.950 7.550 ;
        RECT 14.180 7.280 14.450 7.550 ;
        RECT 27.680 7.280 27.950 7.550 ;
        RECT 41.180 7.280 41.450 7.550 ;
        RECT 54.680 7.280 54.950 7.550 ;
        RECT 68.180 7.280 68.450 7.550 ;
        RECT 81.680 7.280 81.950 7.550 ;
        RECT 95.180 7.280 95.450 7.550 ;
        RECT 108.680 7.280 108.950 7.550 ;
        RECT 122.180 7.280 122.450 7.550 ;
        RECT 135.680 7.280 135.950 7.550 ;
        RECT 149.180 7.280 149.450 7.550 ;
        RECT 162.680 7.280 162.950 7.550 ;
        RECT 176.180 7.280 176.450 7.550 ;
        RECT 189.680 7.280 189.950 7.550 ;
        RECT 203.180 7.280 203.450 7.550 ;
        RECT 216.680 7.280 216.950 7.550 ;
        RECT 7.440 6.380 7.690 6.630 ;
        RECT 20.940 6.380 21.190 6.630 ;
        RECT 34.440 6.380 34.690 6.630 ;
        RECT 47.940 6.380 48.190 6.630 ;
        RECT 61.440 6.380 61.690 6.630 ;
        RECT 74.940 6.380 75.190 6.630 ;
        RECT 88.440 6.380 88.690 6.630 ;
        RECT 101.940 6.380 102.190 6.630 ;
        RECT 115.440 6.380 115.690 6.630 ;
        RECT 128.940 6.380 129.190 6.630 ;
        RECT 142.440 6.380 142.690 6.630 ;
        RECT 155.940 6.380 156.190 6.630 ;
        RECT 169.440 6.380 169.690 6.630 ;
        RECT 182.940 6.380 183.190 6.630 ;
        RECT 196.440 6.380 196.690 6.630 ;
        RECT 209.940 6.380 210.190 6.630 ;
      LAYER met1 ;
        RECT 0.580 7.200 1.040 7.640 ;
        RECT 0.580 7.190 1.050 7.200 ;
        RECT 0.590 6.720 1.050 7.190 ;
        RECT 7.330 6.270 7.800 7.200 ;
        RECT 14.080 6.720 14.550 7.640 ;
        RECT 20.830 6.270 21.300 7.200 ;
        RECT 27.580 6.720 28.050 7.640 ;
        RECT 34.330 6.270 34.800 7.200 ;
        RECT 41.080 6.720 41.550 7.640 ;
        RECT 47.830 6.270 48.300 7.200 ;
        RECT 54.580 6.720 55.050 7.640 ;
        RECT 61.330 6.270 61.800 7.200 ;
        RECT 68.080 6.720 68.550 7.640 ;
        RECT 74.830 6.270 75.300 7.200 ;
        RECT 81.580 6.720 82.050 7.640 ;
        RECT 88.330 6.270 88.800 7.200 ;
        RECT 95.080 6.720 95.550 7.640 ;
        RECT 101.830 6.270 102.300 7.200 ;
        RECT 108.580 6.720 109.050 7.640 ;
        RECT 115.330 6.270 115.800 7.200 ;
        RECT 122.080 6.720 122.550 7.640 ;
        RECT 128.830 6.270 129.300 7.200 ;
        RECT 135.580 6.720 136.050 7.640 ;
        RECT 142.330 6.270 142.800 7.200 ;
        RECT 149.080 6.720 149.550 7.640 ;
        RECT 155.830 6.270 156.300 7.200 ;
        RECT 162.580 6.720 163.050 7.640 ;
        RECT 169.330 6.270 169.800 7.200 ;
        RECT 176.080 6.720 176.550 7.640 ;
        RECT 182.830 6.270 183.300 7.200 ;
        RECT 189.580 6.720 190.050 7.640 ;
        RECT 196.330 6.270 196.800 7.200 ;
        RECT 203.080 6.720 203.550 7.640 ;
        RECT 216.590 7.200 217.050 7.640 ;
        RECT 209.830 6.270 210.300 7.200 ;
        RECT 216.580 7.190 217.050 7.200 ;
        RECT 216.580 6.720 217.040 7.190 ;
      LAYER via ;
        RECT 0.680 6.780 0.950 7.050 ;
        RECT 7.430 6.800 7.700 7.070 ;
        RECT 14.180 6.780 14.450 7.050 ;
        RECT 20.930 6.830 21.200 7.100 ;
        RECT 27.680 6.780 27.950 7.050 ;
        RECT 34.430 6.830 34.700 7.100 ;
        RECT 41.180 6.780 41.450 7.050 ;
        RECT 47.930 6.800 48.200 7.070 ;
        RECT 54.680 6.780 54.950 7.050 ;
        RECT 61.430 6.800 61.700 7.070 ;
        RECT 68.180 6.780 68.450 7.050 ;
        RECT 74.930 6.830 75.200 7.100 ;
        RECT 81.680 6.780 81.950 7.050 ;
        RECT 88.430 6.830 88.700 7.100 ;
        RECT 95.180 6.780 95.450 7.050 ;
        RECT 101.930 6.800 102.200 7.070 ;
        RECT 108.680 6.780 108.950 7.050 ;
        RECT 115.430 6.800 115.700 7.070 ;
        RECT 122.180 6.780 122.450 7.050 ;
        RECT 128.930 6.830 129.200 7.100 ;
        RECT 135.680 6.780 135.950 7.050 ;
        RECT 142.430 6.830 142.700 7.100 ;
        RECT 149.180 6.780 149.450 7.050 ;
        RECT 155.930 6.800 156.200 7.070 ;
        RECT 162.680 6.780 162.950 7.050 ;
        RECT 169.430 6.800 169.700 7.070 ;
        RECT 176.180 6.780 176.450 7.050 ;
        RECT 182.930 6.830 183.200 7.100 ;
        RECT 189.680 6.780 189.950 7.050 ;
        RECT 196.430 6.830 196.700 7.100 ;
        RECT 203.180 6.780 203.450 7.050 ;
        RECT 209.930 6.800 210.200 7.070 ;
        RECT 216.680 6.780 216.950 7.050 ;
      LAYER met2 ;
        RECT 0.880 7.200 1.250 7.210 ;
        RECT 14.040 7.200 41.590 7.210 ;
        RECT 68.040 7.200 95.590 7.210 ;
        RECT 122.040 7.200 149.590 7.210 ;
        RECT 176.040 7.200 203.590 7.210 ;
        RECT 0.590 7.190 217.040 7.200 ;
        RECT 0.580 6.690 217.050 7.190 ;
        RECT 0.580 6.680 14.590 6.690 ;
        RECT 41.040 6.680 68.590 6.690 ;
        RECT 95.040 6.680 122.590 6.690 ;
        RECT 149.040 6.680 176.590 6.690 ;
        RECT 203.040 6.680 217.050 6.690 ;
        RECT 0.580 6.670 1.060 6.680 ;
        RECT 108.570 6.670 109.060 6.680 ;
        RECT 216.570 6.670 217.050 6.680 ;
    END
  END WL5
  PIN WL6
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER li1 ;
        RECT 7.340 5.390 7.790 5.840 ;
        RECT 20.840 5.390 21.290 5.840 ;
        RECT 34.340 5.390 34.790 5.840 ;
        RECT 47.840 5.390 48.290 5.840 ;
        RECT 61.340 5.390 61.790 5.840 ;
        RECT 74.840 5.390 75.290 5.840 ;
        RECT 88.340 5.390 88.790 5.840 ;
        RECT 101.840 5.390 102.290 5.840 ;
        RECT 115.340 5.390 115.790 5.840 ;
        RECT 128.840 5.390 129.290 5.840 ;
        RECT 142.340 5.390 142.790 5.840 ;
        RECT 155.840 5.390 156.290 5.840 ;
        RECT 169.340 5.390 169.790 5.840 ;
        RECT 182.840 5.390 183.290 5.840 ;
        RECT 196.340 5.390 196.790 5.840 ;
        RECT 209.840 5.390 210.290 5.840 ;
        RECT 0.590 4.480 1.040 4.920 ;
        RECT 14.090 4.480 14.540 4.920 ;
        RECT 27.590 4.480 28.040 4.920 ;
        RECT 41.090 4.480 41.540 4.920 ;
        RECT 54.590 4.480 55.040 4.920 ;
        RECT 68.090 4.480 68.540 4.920 ;
        RECT 81.590 4.480 82.040 4.920 ;
        RECT 95.090 4.480 95.540 4.920 ;
        RECT 108.590 4.480 109.040 4.920 ;
        RECT 122.090 4.480 122.540 4.920 ;
        RECT 135.590 4.480 136.040 4.920 ;
        RECT 149.090 4.480 149.540 4.920 ;
        RECT 162.590 4.480 163.040 4.920 ;
        RECT 176.090 4.480 176.540 4.920 ;
        RECT 189.590 4.480 190.040 4.920 ;
        RECT 203.090 4.480 203.540 4.920 ;
        RECT 216.590 4.480 217.040 4.920 ;
      LAYER mcon ;
        RECT 7.440 5.490 7.690 5.740 ;
        RECT 20.940 5.490 21.190 5.740 ;
        RECT 34.440 5.490 34.690 5.740 ;
        RECT 47.940 5.490 48.190 5.740 ;
        RECT 61.440 5.490 61.690 5.740 ;
        RECT 74.940 5.490 75.190 5.740 ;
        RECT 88.440 5.490 88.690 5.740 ;
        RECT 101.940 5.490 102.190 5.740 ;
        RECT 115.440 5.490 115.690 5.740 ;
        RECT 128.940 5.490 129.190 5.740 ;
        RECT 142.440 5.490 142.690 5.740 ;
        RECT 155.940 5.490 156.190 5.740 ;
        RECT 169.440 5.490 169.690 5.740 ;
        RECT 182.940 5.490 183.190 5.740 ;
        RECT 196.440 5.490 196.690 5.740 ;
        RECT 209.940 5.490 210.190 5.740 ;
        RECT 0.680 4.570 0.950 4.840 ;
        RECT 14.180 4.570 14.450 4.840 ;
        RECT 27.680 4.570 27.950 4.840 ;
        RECT 41.180 4.570 41.450 4.840 ;
        RECT 54.680 4.570 54.950 4.840 ;
        RECT 68.180 4.570 68.450 4.840 ;
        RECT 81.680 4.570 81.950 4.840 ;
        RECT 95.180 4.570 95.450 4.840 ;
        RECT 108.680 4.570 108.950 4.840 ;
        RECT 122.180 4.570 122.450 4.840 ;
        RECT 135.680 4.570 135.950 4.840 ;
        RECT 149.180 4.570 149.450 4.840 ;
        RECT 162.680 4.570 162.950 4.840 ;
        RECT 176.180 4.570 176.450 4.840 ;
        RECT 189.680 4.570 189.950 4.840 ;
        RECT 203.180 4.570 203.450 4.840 ;
        RECT 216.680 4.570 216.950 4.840 ;
      LAYER met1 ;
        RECT 0.590 4.930 1.050 5.400 ;
        RECT 0.580 4.920 1.050 4.930 ;
        RECT 7.330 4.920 7.800 5.850 ;
        RECT 0.580 4.480 1.040 4.920 ;
        RECT 14.080 4.480 14.550 5.400 ;
        RECT 20.830 4.920 21.300 5.850 ;
        RECT 27.580 4.480 28.050 5.400 ;
        RECT 34.330 4.920 34.800 5.850 ;
        RECT 41.080 4.480 41.550 5.400 ;
        RECT 47.830 4.920 48.300 5.850 ;
        RECT 54.580 4.480 55.050 5.400 ;
        RECT 61.330 4.920 61.800 5.850 ;
        RECT 68.080 4.480 68.550 5.400 ;
        RECT 74.830 4.920 75.300 5.850 ;
        RECT 81.580 4.480 82.050 5.400 ;
        RECT 88.330 4.920 88.800 5.850 ;
        RECT 95.080 4.480 95.550 5.400 ;
        RECT 101.830 4.920 102.300 5.850 ;
        RECT 108.580 4.480 109.050 5.400 ;
        RECT 115.330 4.920 115.800 5.850 ;
        RECT 122.080 4.480 122.550 5.400 ;
        RECT 128.830 4.920 129.300 5.850 ;
        RECT 135.580 4.480 136.050 5.400 ;
        RECT 142.330 4.920 142.800 5.850 ;
        RECT 149.080 4.480 149.550 5.400 ;
        RECT 155.830 4.920 156.300 5.850 ;
        RECT 162.580 4.480 163.050 5.400 ;
        RECT 169.330 4.920 169.800 5.850 ;
        RECT 176.080 4.480 176.550 5.400 ;
        RECT 182.830 4.920 183.300 5.850 ;
        RECT 189.580 4.480 190.050 5.400 ;
        RECT 196.330 4.920 196.800 5.850 ;
        RECT 203.080 4.480 203.550 5.400 ;
        RECT 209.830 4.920 210.300 5.850 ;
        RECT 216.580 4.930 217.040 5.400 ;
        RECT 216.580 4.920 217.050 4.930 ;
        RECT 216.590 4.480 217.050 4.920 ;
      LAYER via ;
        RECT 0.680 5.070 0.950 5.340 ;
        RECT 7.430 5.020 7.700 5.290 ;
        RECT 14.180 5.070 14.450 5.340 ;
        RECT 20.930 5.020 21.200 5.290 ;
        RECT 27.680 5.070 27.950 5.340 ;
        RECT 34.430 5.020 34.700 5.290 ;
        RECT 41.180 5.070 41.450 5.340 ;
        RECT 47.930 5.020 48.200 5.290 ;
        RECT 54.680 5.070 54.950 5.340 ;
        RECT 61.430 5.020 61.700 5.290 ;
        RECT 68.180 5.070 68.450 5.340 ;
        RECT 74.930 5.020 75.200 5.290 ;
        RECT 81.680 5.070 81.950 5.340 ;
        RECT 88.430 5.020 88.700 5.290 ;
        RECT 95.180 5.070 95.450 5.340 ;
        RECT 101.930 5.020 102.200 5.290 ;
        RECT 108.680 5.070 108.950 5.340 ;
        RECT 115.430 5.020 115.700 5.290 ;
        RECT 122.180 5.070 122.450 5.340 ;
        RECT 128.930 5.020 129.200 5.290 ;
        RECT 135.680 5.070 135.950 5.340 ;
        RECT 142.430 5.020 142.700 5.290 ;
        RECT 149.180 5.070 149.450 5.340 ;
        RECT 155.930 5.020 156.200 5.290 ;
        RECT 162.680 5.070 162.950 5.340 ;
        RECT 169.430 5.020 169.700 5.290 ;
        RECT 176.180 5.070 176.450 5.340 ;
        RECT 182.930 5.020 183.200 5.290 ;
        RECT 189.680 5.070 189.950 5.340 ;
        RECT 196.430 5.020 196.700 5.290 ;
        RECT 203.180 5.070 203.450 5.340 ;
        RECT 209.930 5.020 210.200 5.290 ;
        RECT 216.680 5.070 216.950 5.340 ;
      LAYER met2 ;
        RECT 0.590 4.910 217.040 5.430 ;
    END
  END WL6
  PIN WL7
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER li1 ;
        RECT 0.590 3.590 1.040 4.030 ;
        RECT 14.090 3.590 14.540 4.030 ;
        RECT 27.590 3.590 28.040 4.030 ;
        RECT 41.090 3.590 41.540 4.030 ;
        RECT 54.590 3.590 55.040 4.030 ;
        RECT 68.090 3.590 68.540 4.030 ;
        RECT 81.590 3.590 82.040 4.030 ;
        RECT 95.090 3.590 95.540 4.030 ;
        RECT 108.590 3.590 109.040 4.030 ;
        RECT 122.090 3.590 122.540 4.030 ;
        RECT 135.590 3.590 136.040 4.030 ;
        RECT 149.090 3.590 149.540 4.030 ;
        RECT 162.590 3.590 163.040 4.030 ;
        RECT 176.090 3.590 176.540 4.030 ;
        RECT 189.590 3.590 190.040 4.030 ;
        RECT 203.090 3.590 203.540 4.030 ;
        RECT 216.590 3.590 217.040 4.030 ;
        RECT 7.340 2.670 7.790 3.120 ;
        RECT 20.840 2.670 21.290 3.120 ;
        RECT 34.340 2.670 34.790 3.120 ;
        RECT 47.840 2.670 48.290 3.120 ;
        RECT 61.340 2.670 61.790 3.120 ;
        RECT 74.840 2.670 75.290 3.120 ;
        RECT 88.340 2.670 88.790 3.120 ;
        RECT 101.840 2.670 102.290 3.120 ;
        RECT 115.340 2.670 115.790 3.120 ;
        RECT 128.840 2.670 129.290 3.120 ;
        RECT 142.340 2.670 142.790 3.120 ;
        RECT 155.840 2.670 156.290 3.120 ;
        RECT 169.340 2.670 169.790 3.120 ;
        RECT 182.840 2.670 183.290 3.120 ;
        RECT 196.340 2.670 196.790 3.120 ;
        RECT 209.840 2.670 210.290 3.120 ;
      LAYER mcon ;
        RECT 0.680 3.670 0.950 3.940 ;
        RECT 14.180 3.670 14.450 3.940 ;
        RECT 27.680 3.670 27.950 3.940 ;
        RECT 41.180 3.670 41.450 3.940 ;
        RECT 54.680 3.670 54.950 3.940 ;
        RECT 68.180 3.670 68.450 3.940 ;
        RECT 81.680 3.670 81.950 3.940 ;
        RECT 95.180 3.670 95.450 3.940 ;
        RECT 108.680 3.670 108.950 3.940 ;
        RECT 122.180 3.670 122.450 3.940 ;
        RECT 135.680 3.670 135.950 3.940 ;
        RECT 149.180 3.670 149.450 3.940 ;
        RECT 162.680 3.670 162.950 3.940 ;
        RECT 176.180 3.670 176.450 3.940 ;
        RECT 189.680 3.670 189.950 3.940 ;
        RECT 203.180 3.670 203.450 3.940 ;
        RECT 216.680 3.670 216.950 3.940 ;
        RECT 7.440 2.770 7.690 3.020 ;
        RECT 20.940 2.770 21.190 3.020 ;
        RECT 34.440 2.770 34.690 3.020 ;
        RECT 47.940 2.770 48.190 3.020 ;
        RECT 61.440 2.770 61.690 3.020 ;
        RECT 74.940 2.770 75.190 3.020 ;
        RECT 88.440 2.770 88.690 3.020 ;
        RECT 101.940 2.770 102.190 3.020 ;
        RECT 115.440 2.770 115.690 3.020 ;
        RECT 128.940 2.770 129.190 3.020 ;
        RECT 142.440 2.770 142.690 3.020 ;
        RECT 155.940 2.770 156.190 3.020 ;
        RECT 169.440 2.770 169.690 3.020 ;
        RECT 182.940 2.770 183.190 3.020 ;
        RECT 196.440 2.770 196.690 3.020 ;
        RECT 209.940 2.770 210.190 3.020 ;
      LAYER met1 ;
        RECT 0.580 3.590 1.040 4.030 ;
        RECT 0.580 3.580 1.050 3.590 ;
        RECT 0.590 3.110 1.050 3.580 ;
        RECT 7.330 2.660 7.800 3.590 ;
        RECT 14.080 3.110 14.550 4.030 ;
        RECT 20.830 2.660 21.300 3.590 ;
        RECT 27.580 3.110 28.050 4.030 ;
        RECT 34.330 2.660 34.800 3.590 ;
        RECT 41.080 3.110 41.550 4.030 ;
        RECT 47.830 2.660 48.300 3.590 ;
        RECT 54.580 3.110 55.050 4.030 ;
        RECT 61.330 2.660 61.800 3.590 ;
        RECT 68.080 3.110 68.550 4.030 ;
        RECT 74.830 2.660 75.300 3.590 ;
        RECT 81.580 3.110 82.050 4.030 ;
        RECT 88.330 2.660 88.800 3.590 ;
        RECT 95.080 3.110 95.550 4.030 ;
        RECT 101.830 2.660 102.300 3.590 ;
        RECT 108.580 3.110 109.050 4.030 ;
        RECT 115.330 2.660 115.800 3.590 ;
        RECT 122.080 3.110 122.550 4.030 ;
        RECT 128.830 2.660 129.300 3.590 ;
        RECT 135.580 3.110 136.050 4.030 ;
        RECT 142.330 2.660 142.800 3.590 ;
        RECT 149.080 3.110 149.550 4.030 ;
        RECT 155.830 2.660 156.300 3.590 ;
        RECT 162.580 3.110 163.050 4.030 ;
        RECT 169.330 2.660 169.800 3.590 ;
        RECT 176.080 3.110 176.550 4.030 ;
        RECT 182.830 2.660 183.300 3.590 ;
        RECT 189.580 3.110 190.050 4.030 ;
        RECT 196.330 2.660 196.800 3.590 ;
        RECT 203.080 3.110 203.550 4.030 ;
        RECT 216.590 3.590 217.050 4.030 ;
        RECT 209.830 2.660 210.300 3.590 ;
        RECT 216.580 3.580 217.050 3.590 ;
        RECT 216.580 3.110 217.040 3.580 ;
      LAYER via ;
        RECT 0.680 3.170 0.950 3.440 ;
        RECT 7.430 3.190 7.700 3.460 ;
        RECT 14.180 3.170 14.450 3.440 ;
        RECT 20.930 3.190 21.200 3.460 ;
        RECT 27.680 3.170 27.950 3.440 ;
        RECT 34.430 3.190 34.700 3.460 ;
        RECT 41.180 3.170 41.450 3.440 ;
        RECT 47.930 3.190 48.200 3.460 ;
        RECT 54.680 3.170 54.950 3.440 ;
        RECT 61.430 3.190 61.700 3.460 ;
        RECT 68.180 3.170 68.450 3.440 ;
        RECT 74.930 3.190 75.200 3.460 ;
        RECT 81.680 3.170 81.950 3.440 ;
        RECT 88.430 3.190 88.700 3.460 ;
        RECT 95.180 3.170 95.450 3.440 ;
        RECT 101.930 3.190 102.200 3.460 ;
        RECT 108.680 3.170 108.950 3.440 ;
        RECT 115.430 3.190 115.700 3.460 ;
        RECT 122.180 3.170 122.450 3.440 ;
        RECT 128.930 3.190 129.200 3.460 ;
        RECT 135.680 3.170 135.950 3.440 ;
        RECT 142.430 3.190 142.700 3.460 ;
        RECT 149.180 3.170 149.450 3.440 ;
        RECT 155.930 3.190 156.200 3.460 ;
        RECT 162.680 3.170 162.950 3.440 ;
        RECT 169.430 3.190 169.700 3.460 ;
        RECT 176.180 3.170 176.450 3.440 ;
        RECT 182.930 3.190 183.200 3.460 ;
        RECT 189.680 3.170 189.950 3.440 ;
        RECT 196.430 3.190 196.700 3.460 ;
        RECT 203.180 3.170 203.450 3.440 ;
        RECT 209.930 3.190 210.200 3.460 ;
        RECT 216.680 3.170 216.950 3.440 ;
      LAYER met2 ;
        RECT 0.590 3.570 217.040 3.590 ;
        RECT 0.580 3.070 217.050 3.570 ;
        RECT 0.580 3.060 1.060 3.070 ;
        RECT 108.570 3.060 109.060 3.070 ;
        RECT 216.570 3.060 217.050 3.070 ;
    END
  END WL7
  PIN WL8
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER li1 ;
        RECT 7.340 1.780 7.790 2.230 ;
        RECT 20.840 1.780 21.290 2.230 ;
        RECT 34.340 1.780 34.790 2.230 ;
        RECT 47.840 1.780 48.290 2.230 ;
        RECT 61.340 1.780 61.790 2.230 ;
        RECT 74.840 1.780 75.290 2.230 ;
        RECT 88.340 1.780 88.790 2.230 ;
        RECT 101.840 1.780 102.290 2.230 ;
        RECT 115.340 1.780 115.790 2.230 ;
        RECT 128.840 1.780 129.290 2.230 ;
        RECT 142.340 1.780 142.790 2.230 ;
        RECT 155.840 1.780 156.290 2.230 ;
        RECT 169.340 1.780 169.790 2.230 ;
        RECT 182.840 1.780 183.290 2.230 ;
        RECT 196.340 1.780 196.790 2.230 ;
        RECT 209.840 1.780 210.290 2.230 ;
        RECT 0.590 0.870 1.040 1.310 ;
        RECT 14.090 0.870 14.540 1.310 ;
        RECT 27.590 0.870 28.040 1.310 ;
        RECT 41.090 0.870 41.540 1.310 ;
        RECT 54.590 0.870 55.040 1.310 ;
        RECT 68.090 0.870 68.540 1.310 ;
        RECT 81.590 0.870 82.040 1.310 ;
        RECT 95.090 0.870 95.540 1.310 ;
        RECT 108.590 0.870 109.040 1.310 ;
        RECT 122.090 0.870 122.540 1.310 ;
        RECT 135.590 0.870 136.040 1.310 ;
        RECT 149.090 0.870 149.540 1.310 ;
        RECT 162.590 0.870 163.040 1.310 ;
        RECT 176.090 0.870 176.540 1.310 ;
        RECT 189.590 0.870 190.040 1.310 ;
        RECT 203.090 0.870 203.540 1.310 ;
        RECT 216.590 0.870 217.040 1.310 ;
      LAYER mcon ;
        RECT 7.440 1.880 7.690 2.130 ;
        RECT 20.940 1.880 21.190 2.130 ;
        RECT 34.440 1.880 34.690 2.130 ;
        RECT 47.940 1.880 48.190 2.130 ;
        RECT 61.440 1.880 61.690 2.130 ;
        RECT 74.940 1.880 75.190 2.130 ;
        RECT 88.440 1.880 88.690 2.130 ;
        RECT 101.940 1.880 102.190 2.130 ;
        RECT 115.440 1.880 115.690 2.130 ;
        RECT 128.940 1.880 129.190 2.130 ;
        RECT 142.440 1.880 142.690 2.130 ;
        RECT 155.940 1.880 156.190 2.130 ;
        RECT 169.440 1.880 169.690 2.130 ;
        RECT 182.940 1.880 183.190 2.130 ;
        RECT 196.440 1.880 196.690 2.130 ;
        RECT 209.940 1.880 210.190 2.130 ;
        RECT 0.680 0.960 0.950 1.230 ;
        RECT 14.180 0.960 14.450 1.230 ;
        RECT 27.680 0.960 27.950 1.230 ;
        RECT 41.180 0.960 41.450 1.230 ;
        RECT 54.680 0.960 54.950 1.230 ;
        RECT 68.180 0.960 68.450 1.230 ;
        RECT 81.680 0.960 81.950 1.230 ;
        RECT 95.180 0.960 95.450 1.230 ;
        RECT 108.680 0.960 108.950 1.230 ;
        RECT 122.180 0.960 122.450 1.230 ;
        RECT 135.680 0.960 135.950 1.230 ;
        RECT 149.180 0.960 149.450 1.230 ;
        RECT 162.680 0.960 162.950 1.230 ;
        RECT 176.180 0.960 176.450 1.230 ;
        RECT 189.680 0.960 189.950 1.230 ;
        RECT 203.180 0.960 203.450 1.230 ;
        RECT 216.680 0.960 216.950 1.230 ;
      LAYER met1 ;
        RECT 0.590 1.320 1.050 1.790 ;
        RECT 0.580 1.310 1.050 1.320 ;
        RECT 7.330 1.310 7.800 2.240 ;
        RECT 0.580 0.870 1.040 1.310 ;
        RECT 14.080 0.870 14.550 1.790 ;
        RECT 20.830 1.310 21.300 2.240 ;
        RECT 27.580 0.870 28.050 1.790 ;
        RECT 34.330 1.310 34.800 2.240 ;
        RECT 41.080 0.870 41.550 1.790 ;
        RECT 47.830 1.310 48.300 2.240 ;
        RECT 54.580 0.870 55.050 1.790 ;
        RECT 61.330 1.310 61.800 2.240 ;
        RECT 68.080 0.870 68.550 1.790 ;
        RECT 74.830 1.310 75.300 2.240 ;
        RECT 81.580 0.870 82.050 1.790 ;
        RECT 88.330 1.310 88.800 2.240 ;
        RECT 95.080 0.870 95.550 1.790 ;
        RECT 101.830 1.310 102.300 2.240 ;
        RECT 108.580 0.870 109.050 1.790 ;
        RECT 115.330 1.310 115.800 2.240 ;
        RECT 122.080 0.870 122.550 1.790 ;
        RECT 128.830 1.310 129.300 2.240 ;
        RECT 135.580 0.870 136.050 1.790 ;
        RECT 142.330 1.310 142.800 2.240 ;
        RECT 149.080 0.870 149.550 1.790 ;
        RECT 155.830 1.310 156.300 2.240 ;
        RECT 162.580 0.870 163.050 1.790 ;
        RECT 169.330 1.310 169.800 2.240 ;
        RECT 176.080 0.870 176.550 1.790 ;
        RECT 182.830 1.310 183.300 2.240 ;
        RECT 189.580 0.870 190.050 1.790 ;
        RECT 196.330 1.310 196.800 2.240 ;
        RECT 203.080 0.870 203.550 1.790 ;
        RECT 209.830 1.310 210.300 2.240 ;
        RECT 216.580 1.320 217.040 1.790 ;
        RECT 216.580 1.310 217.050 1.320 ;
        RECT 216.590 0.870 217.050 1.310 ;
      LAYER via ;
        RECT 0.680 1.460 0.950 1.730 ;
        RECT 7.430 1.440 7.700 1.710 ;
        RECT 14.180 1.460 14.450 1.730 ;
        RECT 20.930 1.440 21.200 1.710 ;
        RECT 27.680 1.460 27.950 1.730 ;
        RECT 34.430 1.440 34.700 1.710 ;
        RECT 41.180 1.460 41.450 1.730 ;
        RECT 47.930 1.440 48.200 1.710 ;
        RECT 54.680 1.460 54.950 1.730 ;
        RECT 61.430 1.440 61.700 1.710 ;
        RECT 68.180 1.460 68.450 1.730 ;
        RECT 74.930 1.440 75.200 1.710 ;
        RECT 81.680 1.460 81.950 1.730 ;
        RECT 88.430 1.440 88.700 1.710 ;
        RECT 95.180 1.460 95.450 1.730 ;
        RECT 101.930 1.440 102.200 1.710 ;
        RECT 108.680 1.460 108.950 1.730 ;
        RECT 115.430 1.440 115.700 1.710 ;
        RECT 122.180 1.460 122.450 1.730 ;
        RECT 128.930 1.440 129.200 1.710 ;
        RECT 135.680 1.460 135.950 1.730 ;
        RECT 142.430 1.440 142.700 1.710 ;
        RECT 149.180 1.460 149.450 1.730 ;
        RECT 155.930 1.440 156.200 1.710 ;
        RECT 162.680 1.460 162.950 1.730 ;
        RECT 169.430 1.440 169.700 1.710 ;
        RECT 176.180 1.460 176.450 1.730 ;
        RECT 182.930 1.440 183.200 1.710 ;
        RECT 189.680 1.460 189.950 1.730 ;
        RECT 196.430 1.440 196.700 1.710 ;
        RECT 203.180 1.460 203.450 1.730 ;
        RECT 209.930 1.440 210.200 1.710 ;
        RECT 216.680 1.460 216.950 1.730 ;
      LAYER met2 ;
        RECT 0.580 1.830 1.060 1.840 ;
        RECT 108.570 1.830 109.060 1.840 ;
        RECT 216.570 1.830 217.050 1.840 ;
        RECT 0.580 1.330 217.050 1.830 ;
        RECT 0.590 1.310 217.040 1.330 ;
    END
  END WL8
  PIN WL9
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER li1 ;
        RECT 0.590 -0.020 1.040 0.420 ;
        RECT 14.090 -0.020 14.540 0.420 ;
        RECT 27.590 -0.020 28.040 0.420 ;
        RECT 41.090 -0.020 41.540 0.420 ;
        RECT 54.590 -0.020 55.040 0.420 ;
        RECT 68.090 -0.020 68.540 0.420 ;
        RECT 81.590 -0.020 82.040 0.420 ;
        RECT 95.090 -0.020 95.540 0.420 ;
        RECT 108.590 -0.020 109.040 0.420 ;
        RECT 122.090 -0.020 122.540 0.420 ;
        RECT 135.590 -0.020 136.040 0.420 ;
        RECT 149.090 -0.020 149.540 0.420 ;
        RECT 162.590 -0.020 163.040 0.420 ;
        RECT 176.090 -0.020 176.540 0.420 ;
        RECT 189.590 -0.020 190.040 0.420 ;
        RECT 203.090 -0.020 203.540 0.420 ;
        RECT 216.590 -0.020 217.040 0.420 ;
        RECT 7.340 -0.940 7.790 -0.490 ;
        RECT 20.840 -0.940 21.290 -0.490 ;
        RECT 34.340 -0.940 34.790 -0.490 ;
        RECT 47.840 -0.940 48.290 -0.490 ;
        RECT 61.340 -0.940 61.790 -0.490 ;
        RECT 74.840 -0.940 75.290 -0.490 ;
        RECT 88.340 -0.940 88.790 -0.490 ;
        RECT 101.840 -0.940 102.290 -0.490 ;
        RECT 115.340 -0.940 115.790 -0.490 ;
        RECT 128.840 -0.940 129.290 -0.490 ;
        RECT 142.340 -0.940 142.790 -0.490 ;
        RECT 155.840 -0.940 156.290 -0.490 ;
        RECT 169.340 -0.940 169.790 -0.490 ;
        RECT 182.840 -0.940 183.290 -0.490 ;
        RECT 196.340 -0.940 196.790 -0.490 ;
        RECT 209.840 -0.940 210.290 -0.490 ;
      LAYER mcon ;
        RECT 0.680 0.060 0.950 0.330 ;
        RECT 14.180 0.060 14.450 0.330 ;
        RECT 27.680 0.060 27.950 0.330 ;
        RECT 41.180 0.060 41.450 0.330 ;
        RECT 54.680 0.060 54.950 0.330 ;
        RECT 68.180 0.060 68.450 0.330 ;
        RECT 81.680 0.060 81.950 0.330 ;
        RECT 95.180 0.060 95.450 0.330 ;
        RECT 108.680 0.060 108.950 0.330 ;
        RECT 122.180 0.060 122.450 0.330 ;
        RECT 135.680 0.060 135.950 0.330 ;
        RECT 149.180 0.060 149.450 0.330 ;
        RECT 162.680 0.060 162.950 0.330 ;
        RECT 176.180 0.060 176.450 0.330 ;
        RECT 189.680 0.060 189.950 0.330 ;
        RECT 203.180 0.060 203.450 0.330 ;
        RECT 216.680 0.060 216.950 0.330 ;
        RECT 7.440 -0.840 7.690 -0.590 ;
        RECT 20.940 -0.840 21.190 -0.590 ;
        RECT 34.440 -0.840 34.690 -0.590 ;
        RECT 47.940 -0.840 48.190 -0.590 ;
        RECT 61.440 -0.840 61.690 -0.590 ;
        RECT 74.940 -0.840 75.190 -0.590 ;
        RECT 88.440 -0.840 88.690 -0.590 ;
        RECT 101.940 -0.840 102.190 -0.590 ;
        RECT 115.440 -0.840 115.690 -0.590 ;
        RECT 128.940 -0.840 129.190 -0.590 ;
        RECT 142.440 -0.840 142.690 -0.590 ;
        RECT 155.940 -0.840 156.190 -0.590 ;
        RECT 169.440 -0.840 169.690 -0.590 ;
        RECT 182.940 -0.840 183.190 -0.590 ;
        RECT 196.440 -0.840 196.690 -0.590 ;
        RECT 209.940 -0.840 210.190 -0.590 ;
      LAYER met1 ;
        RECT 0.580 -0.020 1.040 0.420 ;
        RECT 0.580 -0.030 1.050 -0.020 ;
        RECT 0.590 -0.500 1.050 -0.030 ;
        RECT 7.330 -0.950 7.800 -0.020 ;
        RECT 14.080 -0.500 14.550 0.420 ;
        RECT 20.830 -0.950 21.300 -0.020 ;
        RECT 27.580 -0.500 28.050 0.420 ;
        RECT 34.330 -0.950 34.800 -0.020 ;
        RECT 41.080 -0.500 41.550 0.420 ;
        RECT 47.830 -0.950 48.300 -0.020 ;
        RECT 54.580 -0.500 55.050 0.420 ;
        RECT 61.330 -0.950 61.800 -0.020 ;
        RECT 68.080 -0.500 68.550 0.420 ;
        RECT 74.830 -0.950 75.300 -0.020 ;
        RECT 81.580 -0.500 82.050 0.420 ;
        RECT 88.330 -0.950 88.800 -0.020 ;
        RECT 95.080 -0.500 95.550 0.420 ;
        RECT 101.830 -0.950 102.300 -0.020 ;
        RECT 108.580 -0.500 109.050 0.420 ;
        RECT 115.330 -0.950 115.800 -0.020 ;
        RECT 122.080 -0.500 122.550 0.420 ;
        RECT 128.830 -0.950 129.300 -0.020 ;
        RECT 135.580 -0.500 136.050 0.420 ;
        RECT 142.330 -0.950 142.800 -0.020 ;
        RECT 149.080 -0.500 149.550 0.420 ;
        RECT 155.830 -0.950 156.300 -0.020 ;
        RECT 162.580 -0.500 163.050 0.420 ;
        RECT 169.330 -0.950 169.800 -0.020 ;
        RECT 176.080 -0.500 176.550 0.420 ;
        RECT 182.830 -0.950 183.300 -0.020 ;
        RECT 189.580 -0.500 190.050 0.420 ;
        RECT 196.330 -0.950 196.800 -0.020 ;
        RECT 203.080 -0.500 203.550 0.420 ;
        RECT 216.590 -0.020 217.050 0.420 ;
        RECT 209.830 -0.950 210.300 -0.020 ;
        RECT 216.580 -0.030 217.050 -0.020 ;
        RECT 216.580 -0.500 217.040 -0.030 ;
      LAYER via ;
        RECT 0.680 -0.440 0.950 -0.170 ;
        RECT 7.430 -0.390 7.700 -0.120 ;
        RECT 14.180 -0.440 14.450 -0.170 ;
        RECT 20.930 -0.390 21.200 -0.120 ;
        RECT 27.680 -0.440 27.950 -0.170 ;
        RECT 34.430 -0.390 34.700 -0.120 ;
        RECT 41.180 -0.440 41.450 -0.170 ;
        RECT 47.930 -0.390 48.200 -0.120 ;
        RECT 54.680 -0.440 54.950 -0.170 ;
        RECT 61.430 -0.390 61.700 -0.120 ;
        RECT 68.180 -0.440 68.450 -0.170 ;
        RECT 74.930 -0.390 75.200 -0.120 ;
        RECT 81.680 -0.440 81.950 -0.170 ;
        RECT 88.430 -0.390 88.700 -0.120 ;
        RECT 95.180 -0.440 95.450 -0.170 ;
        RECT 101.930 -0.390 102.200 -0.120 ;
        RECT 108.680 -0.440 108.950 -0.170 ;
        RECT 115.430 -0.390 115.700 -0.120 ;
        RECT 122.180 -0.440 122.450 -0.170 ;
        RECT 128.930 -0.390 129.200 -0.120 ;
        RECT 135.680 -0.440 135.950 -0.170 ;
        RECT 142.430 -0.390 142.700 -0.120 ;
        RECT 149.180 -0.440 149.450 -0.170 ;
        RECT 155.930 -0.390 156.200 -0.120 ;
        RECT 162.680 -0.440 162.950 -0.170 ;
        RECT 169.430 -0.390 169.700 -0.120 ;
        RECT 176.180 -0.440 176.450 -0.170 ;
        RECT 182.930 -0.390 183.200 -0.120 ;
        RECT 189.680 -0.440 189.950 -0.170 ;
        RECT 196.430 -0.390 196.700 -0.120 ;
        RECT 203.180 -0.440 203.450 -0.170 ;
        RECT 209.930 -0.390 210.200 -0.120 ;
        RECT 216.680 -0.440 216.950 -0.170 ;
      LAYER met2 ;
        RECT 0.590 -0.530 217.040 -0.010 ;
    END
  END WL9
  PIN WL10
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER li1 ;
        RECT 7.340 -1.830 7.790 -1.380 ;
        RECT 20.840 -1.830 21.290 -1.380 ;
        RECT 34.340 -1.830 34.790 -1.380 ;
        RECT 47.840 -1.830 48.290 -1.380 ;
        RECT 61.340 -1.830 61.790 -1.380 ;
        RECT 74.840 -1.830 75.290 -1.380 ;
        RECT 88.340 -1.830 88.790 -1.380 ;
        RECT 101.840 -1.830 102.290 -1.380 ;
        RECT 115.340 -1.830 115.790 -1.380 ;
        RECT 128.840 -1.830 129.290 -1.380 ;
        RECT 142.340 -1.830 142.790 -1.380 ;
        RECT 155.840 -1.830 156.290 -1.380 ;
        RECT 169.340 -1.830 169.790 -1.380 ;
        RECT 182.840 -1.830 183.290 -1.380 ;
        RECT 196.340 -1.830 196.790 -1.380 ;
        RECT 209.840 -1.830 210.290 -1.380 ;
        RECT 0.590 -2.740 1.040 -2.300 ;
        RECT 14.090 -2.740 14.540 -2.300 ;
        RECT 27.590 -2.740 28.040 -2.300 ;
        RECT 41.090 -2.740 41.540 -2.300 ;
        RECT 54.590 -2.740 55.040 -2.300 ;
        RECT 68.090 -2.740 68.540 -2.300 ;
        RECT 81.590 -2.740 82.040 -2.300 ;
        RECT 95.090 -2.740 95.540 -2.300 ;
        RECT 108.590 -2.740 109.040 -2.300 ;
        RECT 122.090 -2.740 122.540 -2.300 ;
        RECT 135.590 -2.740 136.040 -2.300 ;
        RECT 149.090 -2.740 149.540 -2.300 ;
        RECT 162.590 -2.740 163.040 -2.300 ;
        RECT 176.090 -2.740 176.540 -2.300 ;
        RECT 189.590 -2.740 190.040 -2.300 ;
        RECT 203.090 -2.740 203.540 -2.300 ;
        RECT 216.590 -2.740 217.040 -2.300 ;
      LAYER mcon ;
        RECT 7.440 -1.730 7.690 -1.480 ;
        RECT 20.940 -1.730 21.190 -1.480 ;
        RECT 34.440 -1.730 34.690 -1.480 ;
        RECT 47.940 -1.730 48.190 -1.480 ;
        RECT 61.440 -1.730 61.690 -1.480 ;
        RECT 74.940 -1.730 75.190 -1.480 ;
        RECT 88.440 -1.730 88.690 -1.480 ;
        RECT 101.940 -1.730 102.190 -1.480 ;
        RECT 115.440 -1.730 115.690 -1.480 ;
        RECT 128.940 -1.730 129.190 -1.480 ;
        RECT 142.440 -1.730 142.690 -1.480 ;
        RECT 155.940 -1.730 156.190 -1.480 ;
        RECT 169.440 -1.730 169.690 -1.480 ;
        RECT 182.940 -1.730 183.190 -1.480 ;
        RECT 196.440 -1.730 196.690 -1.480 ;
        RECT 209.940 -1.730 210.190 -1.480 ;
        RECT 0.680 -2.650 0.950 -2.380 ;
        RECT 14.180 -2.650 14.450 -2.380 ;
        RECT 27.680 -2.650 27.950 -2.380 ;
        RECT 41.180 -2.650 41.450 -2.380 ;
        RECT 54.680 -2.650 54.950 -2.380 ;
        RECT 68.180 -2.650 68.450 -2.380 ;
        RECT 81.680 -2.650 81.950 -2.380 ;
        RECT 95.180 -2.650 95.450 -2.380 ;
        RECT 108.680 -2.650 108.950 -2.380 ;
        RECT 122.180 -2.650 122.450 -2.380 ;
        RECT 135.680 -2.650 135.950 -2.380 ;
        RECT 149.180 -2.650 149.450 -2.380 ;
        RECT 162.680 -2.650 162.950 -2.380 ;
        RECT 176.180 -2.650 176.450 -2.380 ;
        RECT 189.680 -2.650 189.950 -2.380 ;
        RECT 203.180 -2.650 203.450 -2.380 ;
        RECT 216.680 -2.650 216.950 -2.380 ;
      LAYER met1 ;
        RECT 0.590 -2.290 1.050 -1.820 ;
        RECT 0.580 -2.300 1.050 -2.290 ;
        RECT 7.330 -2.300 7.800 -1.370 ;
        RECT 0.580 -2.740 1.040 -2.300 ;
        RECT 14.080 -2.740 14.550 -1.820 ;
        RECT 20.830 -2.300 21.300 -1.370 ;
        RECT 27.580 -2.740 28.050 -1.820 ;
        RECT 34.330 -2.300 34.800 -1.370 ;
        RECT 41.080 -2.740 41.550 -1.820 ;
        RECT 47.830 -2.300 48.300 -1.370 ;
        RECT 54.580 -2.740 55.050 -1.820 ;
        RECT 61.330 -2.300 61.800 -1.370 ;
        RECT 68.080 -2.740 68.550 -1.820 ;
        RECT 74.830 -2.300 75.300 -1.370 ;
        RECT 81.580 -2.740 82.050 -1.820 ;
        RECT 88.330 -2.300 88.800 -1.370 ;
        RECT 95.080 -2.740 95.550 -1.820 ;
        RECT 101.830 -2.300 102.300 -1.370 ;
        RECT 108.580 -2.740 109.050 -1.820 ;
        RECT 115.330 -2.300 115.800 -1.370 ;
        RECT 122.080 -2.740 122.550 -1.820 ;
        RECT 128.830 -2.300 129.300 -1.370 ;
        RECT 135.580 -2.740 136.050 -1.820 ;
        RECT 142.330 -2.300 142.800 -1.370 ;
        RECT 149.080 -2.740 149.550 -1.820 ;
        RECT 155.830 -2.300 156.300 -1.370 ;
        RECT 162.580 -2.740 163.050 -1.820 ;
        RECT 169.330 -2.300 169.800 -1.370 ;
        RECT 176.080 -2.740 176.550 -1.820 ;
        RECT 182.830 -2.300 183.300 -1.370 ;
        RECT 189.580 -2.740 190.050 -1.820 ;
        RECT 196.330 -2.300 196.800 -1.370 ;
        RECT 203.080 -2.740 203.550 -1.820 ;
        RECT 209.830 -2.300 210.300 -1.370 ;
        RECT 216.580 -2.290 217.040 -1.820 ;
        RECT 216.580 -2.300 217.050 -2.290 ;
        RECT 216.590 -2.740 217.050 -2.300 ;
      LAYER via ;
        RECT 0.680 -2.150 0.950 -1.880 ;
        RECT 7.430 -2.170 7.700 -1.900 ;
        RECT 14.180 -2.150 14.450 -1.880 ;
        RECT 20.930 -2.200 21.200 -1.930 ;
        RECT 27.680 -2.150 27.950 -1.880 ;
        RECT 34.430 -2.200 34.700 -1.930 ;
        RECT 41.180 -2.150 41.450 -1.880 ;
        RECT 47.930 -2.170 48.200 -1.900 ;
        RECT 54.680 -2.150 54.950 -1.880 ;
        RECT 61.430 -2.170 61.700 -1.900 ;
        RECT 68.180 -2.150 68.450 -1.880 ;
        RECT 74.930 -2.200 75.200 -1.930 ;
        RECT 81.680 -2.150 81.950 -1.880 ;
        RECT 88.430 -2.200 88.700 -1.930 ;
        RECT 95.180 -2.150 95.450 -1.880 ;
        RECT 101.930 -2.170 102.200 -1.900 ;
        RECT 108.680 -2.150 108.950 -1.880 ;
        RECT 115.430 -2.170 115.700 -1.900 ;
        RECT 122.180 -2.150 122.450 -1.880 ;
        RECT 128.930 -2.200 129.200 -1.930 ;
        RECT 135.680 -2.150 135.950 -1.880 ;
        RECT 142.430 -2.200 142.700 -1.930 ;
        RECT 149.180 -2.150 149.450 -1.880 ;
        RECT 155.930 -2.170 156.200 -1.900 ;
        RECT 162.680 -2.150 162.950 -1.880 ;
        RECT 169.430 -2.170 169.700 -1.900 ;
        RECT 176.180 -2.150 176.450 -1.880 ;
        RECT 182.930 -2.200 183.200 -1.930 ;
        RECT 189.680 -2.150 189.950 -1.880 ;
        RECT 196.430 -2.200 196.700 -1.930 ;
        RECT 203.180 -2.150 203.450 -1.880 ;
        RECT 209.930 -2.170 210.200 -1.900 ;
        RECT 216.680 -2.150 216.950 -1.880 ;
      LAYER met2 ;
        RECT 0.580 -1.780 1.060 -1.770 ;
        RECT 108.570 -1.780 109.060 -1.770 ;
        RECT 216.570 -1.780 217.050 -1.770 ;
        RECT 0.580 -1.790 14.590 -1.780 ;
        RECT 41.040 -1.790 68.590 -1.780 ;
        RECT 95.040 -1.790 122.590 -1.780 ;
        RECT 149.040 -1.790 176.590 -1.780 ;
        RECT 203.040 -1.790 217.050 -1.780 ;
        RECT 0.580 -2.290 217.050 -1.790 ;
        RECT 0.590 -2.300 217.040 -2.290 ;
        RECT 14.040 -2.310 41.590 -2.300 ;
        RECT 68.040 -2.310 95.590 -2.300 ;
        RECT 122.040 -2.310 149.590 -2.300 ;
        RECT 176.040 -2.310 203.590 -2.300 ;
    END
  END WL10
  PIN WL11
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER li1 ;
        RECT 0.590 -3.630 1.040 -3.190 ;
        RECT 14.090 -3.630 14.540 -3.190 ;
        RECT 27.590 -3.630 28.040 -3.190 ;
        RECT 41.090 -3.630 41.540 -3.190 ;
        RECT 54.590 -3.630 55.040 -3.190 ;
        RECT 68.090 -3.630 68.540 -3.190 ;
        RECT 81.590 -3.630 82.040 -3.190 ;
        RECT 95.090 -3.630 95.540 -3.190 ;
        RECT 108.590 -3.630 109.040 -3.190 ;
        RECT 122.090 -3.630 122.540 -3.190 ;
        RECT 135.590 -3.630 136.040 -3.190 ;
        RECT 149.090 -3.630 149.540 -3.190 ;
        RECT 162.590 -3.630 163.040 -3.190 ;
        RECT 176.090 -3.630 176.540 -3.190 ;
        RECT 189.590 -3.630 190.040 -3.190 ;
        RECT 203.090 -3.630 203.540 -3.190 ;
        RECT 216.590 -3.630 217.040 -3.190 ;
        RECT 7.340 -4.550 7.790 -4.100 ;
        RECT 20.840 -4.550 21.290 -4.100 ;
        RECT 34.340 -4.550 34.790 -4.100 ;
        RECT 47.840 -4.550 48.290 -4.100 ;
        RECT 61.340 -4.550 61.790 -4.100 ;
        RECT 74.840 -4.550 75.290 -4.100 ;
        RECT 88.340 -4.550 88.790 -4.100 ;
        RECT 101.840 -4.550 102.290 -4.100 ;
        RECT 115.340 -4.550 115.790 -4.100 ;
        RECT 128.840 -4.550 129.290 -4.100 ;
        RECT 142.340 -4.550 142.790 -4.100 ;
        RECT 155.840 -4.550 156.290 -4.100 ;
        RECT 169.340 -4.550 169.790 -4.100 ;
        RECT 182.840 -4.550 183.290 -4.100 ;
        RECT 196.340 -4.550 196.790 -4.100 ;
        RECT 209.840 -4.550 210.290 -4.100 ;
      LAYER mcon ;
        RECT 0.680 -3.550 0.950 -3.280 ;
        RECT 14.180 -3.550 14.450 -3.280 ;
        RECT 27.680 -3.550 27.950 -3.280 ;
        RECT 41.180 -3.550 41.450 -3.280 ;
        RECT 54.680 -3.550 54.950 -3.280 ;
        RECT 68.180 -3.550 68.450 -3.280 ;
        RECT 81.680 -3.550 81.950 -3.280 ;
        RECT 95.180 -3.550 95.450 -3.280 ;
        RECT 108.680 -3.550 108.950 -3.280 ;
        RECT 122.180 -3.550 122.450 -3.280 ;
        RECT 135.680 -3.550 135.950 -3.280 ;
        RECT 149.180 -3.550 149.450 -3.280 ;
        RECT 162.680 -3.550 162.950 -3.280 ;
        RECT 176.180 -3.550 176.450 -3.280 ;
        RECT 189.680 -3.550 189.950 -3.280 ;
        RECT 203.180 -3.550 203.450 -3.280 ;
        RECT 216.680 -3.550 216.950 -3.280 ;
        RECT 7.440 -4.450 7.690 -4.200 ;
        RECT 20.940 -4.450 21.190 -4.200 ;
        RECT 34.440 -4.450 34.690 -4.200 ;
        RECT 47.940 -4.450 48.190 -4.200 ;
        RECT 61.440 -4.450 61.690 -4.200 ;
        RECT 74.940 -4.450 75.190 -4.200 ;
        RECT 88.440 -4.450 88.690 -4.200 ;
        RECT 101.940 -4.450 102.190 -4.200 ;
        RECT 115.440 -4.450 115.690 -4.200 ;
        RECT 128.940 -4.450 129.190 -4.200 ;
        RECT 142.440 -4.450 142.690 -4.200 ;
        RECT 155.940 -4.450 156.190 -4.200 ;
        RECT 169.440 -4.450 169.690 -4.200 ;
        RECT 182.940 -4.450 183.190 -4.200 ;
        RECT 196.440 -4.450 196.690 -4.200 ;
        RECT 209.940 -4.450 210.190 -4.200 ;
      LAYER met1 ;
        RECT 0.580 -3.630 1.040 -3.190 ;
        RECT 0.580 -3.640 1.050 -3.630 ;
        RECT 0.590 -4.110 1.050 -3.640 ;
        RECT 7.330 -4.560 7.800 -3.630 ;
        RECT 14.080 -4.110 14.550 -3.190 ;
        RECT 20.830 -4.560 21.300 -3.630 ;
        RECT 27.580 -4.110 28.050 -3.190 ;
        RECT 34.330 -4.560 34.800 -3.630 ;
        RECT 41.080 -4.110 41.550 -3.190 ;
        RECT 47.830 -4.560 48.300 -3.630 ;
        RECT 54.580 -4.110 55.050 -3.190 ;
        RECT 61.330 -4.560 61.800 -3.630 ;
        RECT 68.080 -4.110 68.550 -3.190 ;
        RECT 74.830 -4.560 75.300 -3.630 ;
        RECT 81.580 -4.110 82.050 -3.190 ;
        RECT 88.330 -4.560 88.800 -3.630 ;
        RECT 95.080 -4.110 95.550 -3.190 ;
        RECT 101.830 -4.560 102.300 -3.630 ;
        RECT 108.580 -4.110 109.050 -3.190 ;
        RECT 115.330 -4.560 115.800 -3.630 ;
        RECT 122.080 -4.110 122.550 -3.190 ;
        RECT 128.830 -4.560 129.300 -3.630 ;
        RECT 135.580 -4.110 136.050 -3.190 ;
        RECT 142.330 -4.560 142.800 -3.630 ;
        RECT 149.080 -4.110 149.550 -3.190 ;
        RECT 155.830 -4.560 156.300 -3.630 ;
        RECT 162.580 -4.110 163.050 -3.190 ;
        RECT 169.330 -4.560 169.800 -3.630 ;
        RECT 176.080 -4.110 176.550 -3.190 ;
        RECT 182.830 -4.560 183.300 -3.630 ;
        RECT 189.580 -4.110 190.050 -3.190 ;
        RECT 196.330 -4.560 196.800 -3.630 ;
        RECT 203.080 -4.110 203.550 -3.190 ;
        RECT 216.590 -3.630 217.050 -3.190 ;
        RECT 209.830 -4.560 210.300 -3.630 ;
        RECT 216.580 -3.640 217.050 -3.630 ;
        RECT 216.580 -4.110 217.040 -3.640 ;
      LAYER via ;
        RECT 0.680 -4.050 0.950 -3.780 ;
        RECT 7.430 -4.000 7.700 -3.730 ;
        RECT 14.180 -4.050 14.450 -3.780 ;
        RECT 20.930 -4.030 21.200 -3.760 ;
        RECT 27.680 -4.050 27.950 -3.780 ;
        RECT 34.430 -4.030 34.700 -3.760 ;
        RECT 41.180 -4.050 41.450 -3.780 ;
        RECT 47.930 -4.000 48.200 -3.730 ;
        RECT 54.680 -4.050 54.950 -3.780 ;
        RECT 61.430 -4.000 61.700 -3.730 ;
        RECT 68.180 -4.050 68.450 -3.780 ;
        RECT 74.930 -4.030 75.200 -3.760 ;
        RECT 81.680 -4.050 81.950 -3.780 ;
        RECT 88.430 -4.030 88.700 -3.760 ;
        RECT 95.180 -4.050 95.450 -3.780 ;
        RECT 101.930 -4.000 102.200 -3.730 ;
        RECT 108.680 -4.050 108.950 -3.780 ;
        RECT 115.430 -4.000 115.700 -3.730 ;
        RECT 122.180 -4.050 122.450 -3.780 ;
        RECT 128.930 -4.030 129.200 -3.760 ;
        RECT 135.680 -4.050 135.950 -3.780 ;
        RECT 142.430 -4.030 142.700 -3.760 ;
        RECT 149.180 -4.050 149.450 -3.780 ;
        RECT 155.930 -4.000 156.200 -3.730 ;
        RECT 162.680 -4.050 162.950 -3.780 ;
        RECT 169.430 -4.000 169.700 -3.730 ;
        RECT 176.180 -4.050 176.450 -3.780 ;
        RECT 182.930 -4.030 183.200 -3.760 ;
        RECT 189.680 -4.050 189.950 -3.780 ;
        RECT 196.430 -4.030 196.700 -3.760 ;
        RECT 203.180 -4.050 203.450 -3.780 ;
        RECT 209.930 -4.000 210.200 -3.730 ;
        RECT 216.680 -4.050 216.950 -3.780 ;
      LAYER met2 ;
        RECT 0.590 -3.630 14.590 -3.620 ;
        RECT 41.040 -3.630 68.590 -3.620 ;
        RECT 95.040 -3.630 122.590 -3.620 ;
        RECT 149.040 -3.630 176.590 -3.620 ;
        RECT 203.040 -3.630 217.040 -3.620 ;
        RECT 0.590 -3.640 217.040 -3.630 ;
        RECT 0.580 -4.140 217.050 -3.640 ;
        RECT 0.580 -4.150 1.060 -4.140 ;
        RECT 14.040 -4.150 41.590 -4.140 ;
        RECT 68.040 -4.150 95.590 -4.140 ;
        RECT 108.570 -4.150 109.060 -4.140 ;
        RECT 122.040 -4.150 149.590 -4.140 ;
        RECT 176.040 -4.150 203.590 -4.140 ;
        RECT 216.570 -4.150 217.050 -4.140 ;
    END
  END WL11
  PIN WL12
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER li1 ;
        RECT 7.340 -5.440 7.790 -4.990 ;
        RECT 20.840 -5.440 21.290 -4.990 ;
        RECT 34.340 -5.440 34.790 -4.990 ;
        RECT 47.840 -5.440 48.290 -4.990 ;
        RECT 61.340 -5.440 61.790 -4.990 ;
        RECT 74.840 -5.440 75.290 -4.990 ;
        RECT 88.340 -5.440 88.790 -4.990 ;
        RECT 101.840 -5.440 102.290 -4.990 ;
        RECT 115.340 -5.440 115.790 -4.990 ;
        RECT 128.840 -5.440 129.290 -4.990 ;
        RECT 142.340 -5.440 142.790 -4.990 ;
        RECT 155.840 -5.440 156.290 -4.990 ;
        RECT 169.340 -5.440 169.790 -4.990 ;
        RECT 182.840 -5.440 183.290 -4.990 ;
        RECT 196.340 -5.440 196.790 -4.990 ;
        RECT 209.840 -5.440 210.290 -4.990 ;
        RECT 0.590 -6.350 1.040 -5.910 ;
        RECT 14.090 -6.350 14.540 -5.910 ;
        RECT 27.590 -6.350 28.040 -5.910 ;
        RECT 41.090 -6.350 41.540 -5.910 ;
        RECT 54.590 -6.350 55.040 -5.910 ;
        RECT 68.090 -6.350 68.540 -5.910 ;
        RECT 81.590 -6.350 82.040 -5.910 ;
        RECT 95.090 -6.350 95.540 -5.910 ;
        RECT 108.590 -6.350 109.040 -5.910 ;
        RECT 122.090 -6.350 122.540 -5.910 ;
        RECT 135.590 -6.350 136.040 -5.910 ;
        RECT 149.090 -6.350 149.540 -5.910 ;
        RECT 162.590 -6.350 163.040 -5.910 ;
        RECT 176.090 -6.350 176.540 -5.910 ;
        RECT 189.590 -6.350 190.040 -5.910 ;
        RECT 203.090 -6.350 203.540 -5.910 ;
        RECT 216.590 -6.350 217.040 -5.910 ;
      LAYER mcon ;
        RECT 7.440 -5.340 7.690 -5.090 ;
        RECT 20.940 -5.340 21.190 -5.090 ;
        RECT 34.440 -5.340 34.690 -5.090 ;
        RECT 47.940 -5.340 48.190 -5.090 ;
        RECT 61.440 -5.340 61.690 -5.090 ;
        RECT 74.940 -5.340 75.190 -5.090 ;
        RECT 88.440 -5.340 88.690 -5.090 ;
        RECT 101.940 -5.340 102.190 -5.090 ;
        RECT 115.440 -5.340 115.690 -5.090 ;
        RECT 128.940 -5.340 129.190 -5.090 ;
        RECT 142.440 -5.340 142.690 -5.090 ;
        RECT 155.940 -5.340 156.190 -5.090 ;
        RECT 169.440 -5.340 169.690 -5.090 ;
        RECT 182.940 -5.340 183.190 -5.090 ;
        RECT 196.440 -5.340 196.690 -5.090 ;
        RECT 209.940 -5.340 210.190 -5.090 ;
        RECT 0.680 -6.260 0.950 -5.990 ;
        RECT 14.180 -6.260 14.450 -5.990 ;
        RECT 27.680 -6.260 27.950 -5.990 ;
        RECT 41.180 -6.260 41.450 -5.990 ;
        RECT 54.680 -6.260 54.950 -5.990 ;
        RECT 68.180 -6.260 68.450 -5.990 ;
        RECT 81.680 -6.260 81.950 -5.990 ;
        RECT 95.180 -6.260 95.450 -5.990 ;
        RECT 108.680 -6.260 108.950 -5.990 ;
        RECT 122.180 -6.260 122.450 -5.990 ;
        RECT 135.680 -6.260 135.950 -5.990 ;
        RECT 149.180 -6.260 149.450 -5.990 ;
        RECT 162.680 -6.260 162.950 -5.990 ;
        RECT 176.180 -6.260 176.450 -5.990 ;
        RECT 189.680 -6.260 189.950 -5.990 ;
        RECT 203.180 -6.260 203.450 -5.990 ;
        RECT 216.680 -6.260 216.950 -5.990 ;
      LAYER met1 ;
        RECT 0.590 -5.900 1.050 -5.430 ;
        RECT 0.580 -5.910 1.050 -5.900 ;
        RECT 7.330 -5.910 7.800 -4.980 ;
        RECT 0.580 -6.350 1.040 -5.910 ;
        RECT 14.080 -6.350 14.550 -5.430 ;
        RECT 20.830 -5.910 21.300 -4.980 ;
        RECT 27.580 -6.350 28.050 -5.430 ;
        RECT 34.330 -5.910 34.800 -4.980 ;
        RECT 41.080 -6.350 41.550 -5.430 ;
        RECT 47.830 -5.910 48.300 -4.980 ;
        RECT 54.580 -6.350 55.050 -5.430 ;
        RECT 61.330 -5.910 61.800 -4.980 ;
        RECT 68.080 -6.350 68.550 -5.430 ;
        RECT 74.830 -5.910 75.300 -4.980 ;
        RECT 81.580 -6.350 82.050 -5.430 ;
        RECT 88.330 -5.910 88.800 -4.980 ;
        RECT 95.080 -6.350 95.550 -5.430 ;
        RECT 101.830 -5.910 102.300 -4.980 ;
        RECT 108.580 -6.350 109.050 -5.430 ;
        RECT 115.330 -5.910 115.800 -4.980 ;
        RECT 122.080 -6.350 122.550 -5.430 ;
        RECT 128.830 -5.910 129.300 -4.980 ;
        RECT 135.580 -6.350 136.050 -5.430 ;
        RECT 142.330 -5.910 142.800 -4.980 ;
        RECT 149.080 -6.350 149.550 -5.430 ;
        RECT 155.830 -5.910 156.300 -4.980 ;
        RECT 162.580 -6.350 163.050 -5.430 ;
        RECT 169.330 -5.910 169.800 -4.980 ;
        RECT 176.080 -6.350 176.550 -5.430 ;
        RECT 182.830 -5.910 183.300 -4.980 ;
        RECT 189.580 -6.350 190.050 -5.430 ;
        RECT 196.330 -5.910 196.800 -4.980 ;
        RECT 203.080 -6.350 203.550 -5.430 ;
        RECT 209.830 -5.910 210.300 -4.980 ;
        RECT 216.580 -5.900 217.040 -5.430 ;
        RECT 216.580 -5.910 217.050 -5.900 ;
        RECT 216.590 -6.350 217.050 -5.910 ;
      LAYER via ;
        RECT 0.680 -5.760 0.950 -5.490 ;
        RECT 7.430 -5.810 7.700 -5.540 ;
        RECT 14.180 -5.760 14.450 -5.490 ;
        RECT 20.930 -5.780 21.200 -5.510 ;
        RECT 27.680 -5.760 27.950 -5.490 ;
        RECT 34.430 -5.780 34.700 -5.510 ;
        RECT 41.180 -5.760 41.450 -5.490 ;
        RECT 47.930 -5.810 48.200 -5.540 ;
        RECT 54.680 -5.760 54.950 -5.490 ;
        RECT 61.430 -5.810 61.700 -5.540 ;
        RECT 68.180 -5.760 68.450 -5.490 ;
        RECT 74.930 -5.780 75.200 -5.510 ;
        RECT 81.680 -5.760 81.950 -5.490 ;
        RECT 88.430 -5.780 88.700 -5.510 ;
        RECT 95.180 -5.760 95.450 -5.490 ;
        RECT 101.930 -5.810 102.200 -5.540 ;
        RECT 108.680 -5.760 108.950 -5.490 ;
        RECT 115.430 -5.810 115.700 -5.540 ;
        RECT 122.180 -5.760 122.450 -5.490 ;
        RECT 128.930 -5.780 129.200 -5.510 ;
        RECT 135.680 -5.760 135.950 -5.490 ;
        RECT 142.430 -5.780 142.700 -5.510 ;
        RECT 149.180 -5.760 149.450 -5.490 ;
        RECT 155.930 -5.810 156.200 -5.540 ;
        RECT 162.680 -5.760 162.950 -5.490 ;
        RECT 169.430 -5.810 169.700 -5.540 ;
        RECT 176.180 -5.760 176.450 -5.490 ;
        RECT 182.930 -5.780 183.200 -5.510 ;
        RECT 189.680 -5.760 189.950 -5.490 ;
        RECT 196.430 -5.780 196.700 -5.510 ;
        RECT 203.180 -5.760 203.450 -5.490 ;
        RECT 209.930 -5.810 210.200 -5.540 ;
        RECT 216.680 -5.760 216.950 -5.490 ;
      LAYER met2 ;
        RECT 0.870 -5.400 1.240 -5.390 ;
        RECT 14.040 -5.400 41.590 -5.390 ;
        RECT 68.040 -5.400 95.590 -5.390 ;
        RECT 122.040 -5.400 149.590 -5.390 ;
        RECT 176.040 -5.400 203.590 -5.390 ;
        RECT 0.590 -5.410 217.040 -5.400 ;
        RECT 0.580 -5.890 217.050 -5.410 ;
        RECT 0.590 -5.910 217.040 -5.890 ;
        RECT 0.590 -5.920 14.590 -5.910 ;
        RECT 41.040 -5.920 68.590 -5.910 ;
        RECT 95.040 -5.920 122.590 -5.910 ;
        RECT 149.040 -5.920 176.590 -5.910 ;
        RECT 203.040 -5.920 217.040 -5.910 ;
    END
  END WL12
  PIN WL13
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER li1 ;
        RECT 0.590 -7.240 1.040 -6.800 ;
        RECT 14.090 -7.240 14.540 -6.800 ;
        RECT 27.590 -7.240 28.040 -6.800 ;
        RECT 41.090 -7.240 41.540 -6.800 ;
        RECT 54.590 -7.240 55.040 -6.800 ;
        RECT 68.090 -7.240 68.540 -6.800 ;
        RECT 81.590 -7.240 82.040 -6.800 ;
        RECT 95.090 -7.240 95.540 -6.800 ;
        RECT 108.590 -7.240 109.040 -6.800 ;
        RECT 122.090 -7.240 122.540 -6.800 ;
        RECT 135.590 -7.240 136.040 -6.800 ;
        RECT 149.090 -7.240 149.540 -6.800 ;
        RECT 162.590 -7.240 163.040 -6.800 ;
        RECT 176.090 -7.240 176.540 -6.800 ;
        RECT 189.590 -7.240 190.040 -6.800 ;
        RECT 203.090 -7.240 203.540 -6.800 ;
        RECT 216.590 -7.240 217.040 -6.800 ;
        RECT 7.340 -8.160 7.790 -7.710 ;
        RECT 20.840 -8.160 21.290 -7.710 ;
        RECT 34.340 -8.160 34.790 -7.710 ;
        RECT 47.840 -8.160 48.290 -7.710 ;
        RECT 61.340 -8.160 61.790 -7.710 ;
        RECT 74.840 -8.160 75.290 -7.710 ;
        RECT 88.340 -8.160 88.790 -7.710 ;
        RECT 101.840 -8.160 102.290 -7.710 ;
        RECT 115.340 -8.160 115.790 -7.710 ;
        RECT 128.840 -8.160 129.290 -7.710 ;
        RECT 142.340 -8.160 142.790 -7.710 ;
        RECT 155.840 -8.160 156.290 -7.710 ;
        RECT 169.340 -8.160 169.790 -7.710 ;
        RECT 182.840 -8.160 183.290 -7.710 ;
        RECT 196.340 -8.160 196.790 -7.710 ;
        RECT 209.840 -8.160 210.290 -7.710 ;
      LAYER mcon ;
        RECT 0.680 -7.160 0.950 -6.890 ;
        RECT 14.180 -7.160 14.450 -6.890 ;
        RECT 27.680 -7.160 27.950 -6.890 ;
        RECT 41.180 -7.160 41.450 -6.890 ;
        RECT 54.680 -7.160 54.950 -6.890 ;
        RECT 68.180 -7.160 68.450 -6.890 ;
        RECT 81.680 -7.160 81.950 -6.890 ;
        RECT 95.180 -7.160 95.450 -6.890 ;
        RECT 108.680 -7.160 108.950 -6.890 ;
        RECT 122.180 -7.160 122.450 -6.890 ;
        RECT 135.680 -7.160 135.950 -6.890 ;
        RECT 149.180 -7.160 149.450 -6.890 ;
        RECT 162.680 -7.160 162.950 -6.890 ;
        RECT 176.180 -7.160 176.450 -6.890 ;
        RECT 189.680 -7.160 189.950 -6.890 ;
        RECT 203.180 -7.160 203.450 -6.890 ;
        RECT 216.680 -7.160 216.950 -6.890 ;
        RECT 7.440 -8.060 7.690 -7.810 ;
        RECT 20.940 -8.060 21.190 -7.810 ;
        RECT 34.440 -8.060 34.690 -7.810 ;
        RECT 47.940 -8.060 48.190 -7.810 ;
        RECT 61.440 -8.060 61.690 -7.810 ;
        RECT 74.940 -8.060 75.190 -7.810 ;
        RECT 88.440 -8.060 88.690 -7.810 ;
        RECT 101.940 -8.060 102.190 -7.810 ;
        RECT 115.440 -8.060 115.690 -7.810 ;
        RECT 128.940 -8.060 129.190 -7.810 ;
        RECT 142.440 -8.060 142.690 -7.810 ;
        RECT 155.940 -8.060 156.190 -7.810 ;
        RECT 169.440 -8.060 169.690 -7.810 ;
        RECT 182.940 -8.060 183.190 -7.810 ;
        RECT 196.440 -8.060 196.690 -7.810 ;
        RECT 209.940 -8.060 210.190 -7.810 ;
      LAYER met1 ;
        RECT 0.580 -7.240 1.040 -6.800 ;
        RECT 0.580 -7.250 1.050 -7.240 ;
        RECT 0.590 -7.720 1.050 -7.250 ;
        RECT 7.330 -8.170 7.800 -7.240 ;
        RECT 14.080 -7.720 14.550 -6.800 ;
        RECT 20.830 -8.170 21.300 -7.240 ;
        RECT 27.580 -7.720 28.050 -6.800 ;
        RECT 34.330 -8.170 34.800 -7.240 ;
        RECT 41.080 -7.720 41.550 -6.800 ;
        RECT 47.830 -8.170 48.300 -7.240 ;
        RECT 54.580 -7.720 55.050 -6.800 ;
        RECT 61.330 -8.170 61.800 -7.240 ;
        RECT 68.080 -7.720 68.550 -6.800 ;
        RECT 74.830 -8.170 75.300 -7.240 ;
        RECT 81.580 -7.720 82.050 -6.800 ;
        RECT 88.330 -8.170 88.800 -7.240 ;
        RECT 95.080 -7.720 95.550 -6.800 ;
        RECT 101.830 -8.170 102.300 -7.240 ;
        RECT 108.580 -7.720 109.050 -6.800 ;
        RECT 115.330 -8.170 115.800 -7.240 ;
        RECT 122.080 -7.720 122.550 -6.800 ;
        RECT 128.830 -8.170 129.300 -7.240 ;
        RECT 135.580 -7.720 136.050 -6.800 ;
        RECT 142.330 -8.170 142.800 -7.240 ;
        RECT 149.080 -7.720 149.550 -6.800 ;
        RECT 155.830 -8.170 156.300 -7.240 ;
        RECT 162.580 -7.720 163.050 -6.800 ;
        RECT 169.330 -8.170 169.800 -7.240 ;
        RECT 176.080 -7.720 176.550 -6.800 ;
        RECT 182.830 -8.170 183.300 -7.240 ;
        RECT 189.580 -7.720 190.050 -6.800 ;
        RECT 196.330 -8.170 196.800 -7.240 ;
        RECT 203.080 -7.720 203.550 -6.800 ;
        RECT 216.590 -7.240 217.050 -6.800 ;
        RECT 209.830 -8.170 210.300 -7.240 ;
        RECT 216.580 -7.250 217.050 -7.240 ;
        RECT 216.580 -7.720 217.040 -7.250 ;
      LAYER via ;
        RECT 0.680 -7.660 0.950 -7.390 ;
        RECT 7.430 -7.640 7.700 -7.370 ;
        RECT 14.180 -7.660 14.450 -7.390 ;
        RECT 20.930 -7.610 21.200 -7.340 ;
        RECT 27.680 -7.660 27.950 -7.390 ;
        RECT 34.430 -7.610 34.700 -7.340 ;
        RECT 41.180 -7.660 41.450 -7.390 ;
        RECT 47.930 -7.640 48.200 -7.370 ;
        RECT 54.680 -7.660 54.950 -7.390 ;
        RECT 61.430 -7.640 61.700 -7.370 ;
        RECT 68.180 -7.660 68.450 -7.390 ;
        RECT 74.930 -7.610 75.200 -7.340 ;
        RECT 81.680 -7.660 81.950 -7.390 ;
        RECT 88.430 -7.610 88.700 -7.340 ;
        RECT 95.180 -7.660 95.450 -7.390 ;
        RECT 101.930 -7.640 102.200 -7.370 ;
        RECT 108.680 -7.660 108.950 -7.390 ;
        RECT 115.430 -7.640 115.700 -7.370 ;
        RECT 122.180 -7.660 122.450 -7.390 ;
        RECT 128.930 -7.610 129.200 -7.340 ;
        RECT 135.680 -7.660 135.950 -7.390 ;
        RECT 142.430 -7.610 142.700 -7.340 ;
        RECT 149.180 -7.660 149.450 -7.390 ;
        RECT 155.930 -7.640 156.200 -7.370 ;
        RECT 162.680 -7.660 162.950 -7.390 ;
        RECT 169.430 -7.640 169.700 -7.370 ;
        RECT 176.180 -7.660 176.450 -7.390 ;
        RECT 182.930 -7.610 183.200 -7.340 ;
        RECT 189.680 -7.660 189.950 -7.390 ;
        RECT 196.430 -7.610 196.700 -7.340 ;
        RECT 203.180 -7.660 203.450 -7.390 ;
        RECT 209.930 -7.640 210.200 -7.370 ;
        RECT 216.680 -7.660 216.950 -7.390 ;
      LAYER met2 ;
        RECT 14.040 -7.240 41.590 -7.230 ;
        RECT 68.040 -7.240 95.590 -7.230 ;
        RECT 122.040 -7.240 149.590 -7.230 ;
        RECT 176.040 -7.240 203.590 -7.230 ;
        RECT 0.590 -7.250 217.040 -7.240 ;
        RECT 0.580 -7.730 217.050 -7.250 ;
        RECT 0.590 -7.750 217.040 -7.730 ;
        RECT 0.590 -7.760 14.590 -7.750 ;
        RECT 41.040 -7.760 68.590 -7.750 ;
        RECT 95.040 -7.760 122.590 -7.750 ;
        RECT 149.040 -7.760 176.590 -7.750 ;
        RECT 203.040 -7.760 217.040 -7.750 ;
        RECT 0.590 -7.770 1.070 -7.760 ;
        RECT 108.560 -7.770 109.070 -7.760 ;
        RECT 216.560 -7.770 217.040 -7.760 ;
    END
  END WL13
  PIN WL14
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER li1 ;
        RECT 7.340 -9.050 7.790 -8.600 ;
        RECT 20.840 -9.050 21.290 -8.600 ;
        RECT 34.340 -9.050 34.790 -8.600 ;
        RECT 47.840 -9.050 48.290 -8.600 ;
        RECT 61.340 -9.050 61.790 -8.600 ;
        RECT 74.840 -9.050 75.290 -8.600 ;
        RECT 88.340 -9.050 88.790 -8.600 ;
        RECT 101.840 -9.050 102.290 -8.600 ;
        RECT 115.340 -9.050 115.790 -8.600 ;
        RECT 128.840 -9.050 129.290 -8.600 ;
        RECT 142.340 -9.050 142.790 -8.600 ;
        RECT 155.840 -9.050 156.290 -8.600 ;
        RECT 169.340 -9.050 169.790 -8.600 ;
        RECT 182.840 -9.050 183.290 -8.600 ;
        RECT 196.340 -9.050 196.790 -8.600 ;
        RECT 209.840 -9.050 210.290 -8.600 ;
        RECT 0.590 -9.960 1.040 -9.520 ;
        RECT 14.090 -9.960 14.540 -9.520 ;
        RECT 27.590 -9.960 28.040 -9.520 ;
        RECT 41.090 -9.960 41.540 -9.520 ;
        RECT 54.590 -9.960 55.040 -9.520 ;
        RECT 68.090 -9.960 68.540 -9.520 ;
        RECT 81.590 -9.960 82.040 -9.520 ;
        RECT 95.090 -9.960 95.540 -9.520 ;
        RECT 108.590 -9.960 109.040 -9.520 ;
        RECT 122.090 -9.960 122.540 -9.520 ;
        RECT 135.590 -9.960 136.040 -9.520 ;
        RECT 149.090 -9.960 149.540 -9.520 ;
        RECT 162.590 -9.960 163.040 -9.520 ;
        RECT 176.090 -9.960 176.540 -9.520 ;
        RECT 189.590 -9.960 190.040 -9.520 ;
        RECT 203.090 -9.960 203.540 -9.520 ;
        RECT 216.590 -9.960 217.040 -9.520 ;
      LAYER mcon ;
        RECT 7.440 -8.950 7.690 -8.700 ;
        RECT 20.940 -8.950 21.190 -8.700 ;
        RECT 34.440 -8.950 34.690 -8.700 ;
        RECT 47.940 -8.950 48.190 -8.700 ;
        RECT 61.440 -8.950 61.690 -8.700 ;
        RECT 74.940 -8.950 75.190 -8.700 ;
        RECT 88.440 -8.950 88.690 -8.700 ;
        RECT 101.940 -8.950 102.190 -8.700 ;
        RECT 115.440 -8.950 115.690 -8.700 ;
        RECT 128.940 -8.950 129.190 -8.700 ;
        RECT 142.440 -8.950 142.690 -8.700 ;
        RECT 155.940 -8.950 156.190 -8.700 ;
        RECT 169.440 -8.950 169.690 -8.700 ;
        RECT 182.940 -8.950 183.190 -8.700 ;
        RECT 196.440 -8.950 196.690 -8.700 ;
        RECT 209.940 -8.950 210.190 -8.700 ;
        RECT 0.680 -9.870 0.950 -9.600 ;
        RECT 14.180 -9.870 14.450 -9.600 ;
        RECT 27.680 -9.870 27.950 -9.600 ;
        RECT 41.180 -9.870 41.450 -9.600 ;
        RECT 54.680 -9.870 54.950 -9.600 ;
        RECT 68.180 -9.870 68.450 -9.600 ;
        RECT 81.680 -9.870 81.950 -9.600 ;
        RECT 95.180 -9.870 95.450 -9.600 ;
        RECT 108.680 -9.870 108.950 -9.600 ;
        RECT 122.180 -9.870 122.450 -9.600 ;
        RECT 135.680 -9.870 135.950 -9.600 ;
        RECT 149.180 -9.870 149.450 -9.600 ;
        RECT 162.680 -9.870 162.950 -9.600 ;
        RECT 176.180 -9.870 176.450 -9.600 ;
        RECT 189.680 -9.870 189.950 -9.600 ;
        RECT 203.180 -9.870 203.450 -9.600 ;
        RECT 216.680 -9.870 216.950 -9.600 ;
      LAYER met1 ;
        RECT 0.590 -9.510 1.050 -9.040 ;
        RECT 0.580 -9.520 1.050 -9.510 ;
        RECT 7.330 -9.520 7.800 -8.590 ;
        RECT 0.580 -9.960 1.040 -9.520 ;
        RECT 14.080 -9.960 14.550 -9.040 ;
        RECT 20.830 -9.520 21.300 -8.590 ;
        RECT 27.580 -9.960 28.050 -9.040 ;
        RECT 34.330 -9.520 34.800 -8.590 ;
        RECT 41.080 -9.960 41.550 -9.040 ;
        RECT 47.830 -9.520 48.300 -8.590 ;
        RECT 54.580 -9.960 55.050 -9.040 ;
        RECT 61.330 -9.520 61.800 -8.590 ;
        RECT 68.080 -9.960 68.550 -9.040 ;
        RECT 74.830 -9.520 75.300 -8.590 ;
        RECT 81.580 -9.960 82.050 -9.040 ;
        RECT 88.330 -9.520 88.800 -8.590 ;
        RECT 95.080 -9.960 95.550 -9.040 ;
        RECT 101.830 -9.520 102.300 -8.590 ;
        RECT 108.580 -9.960 109.050 -9.040 ;
        RECT 115.330 -9.520 115.800 -8.590 ;
        RECT 122.080 -9.960 122.550 -9.040 ;
        RECT 128.830 -9.520 129.300 -8.590 ;
        RECT 135.580 -9.960 136.050 -9.040 ;
        RECT 142.330 -9.520 142.800 -8.590 ;
        RECT 149.080 -9.960 149.550 -9.040 ;
        RECT 155.830 -9.520 156.300 -8.590 ;
        RECT 162.580 -9.960 163.050 -9.040 ;
        RECT 169.330 -9.520 169.800 -8.590 ;
        RECT 176.080 -9.960 176.550 -9.040 ;
        RECT 182.830 -9.520 183.300 -8.590 ;
        RECT 189.580 -9.960 190.050 -9.040 ;
        RECT 196.330 -9.520 196.800 -8.590 ;
        RECT 203.080 -9.960 203.550 -9.040 ;
        RECT 209.830 -9.520 210.300 -8.590 ;
        RECT 216.580 -9.510 217.040 -9.040 ;
        RECT 216.580 -9.520 217.050 -9.510 ;
        RECT 216.590 -9.960 217.050 -9.520 ;
      LAYER via ;
        RECT 0.680 -9.370 0.950 -9.100 ;
        RECT 7.430 -9.420 7.700 -9.150 ;
        RECT 14.180 -9.370 14.450 -9.100 ;
        RECT 20.930 -9.420 21.200 -9.150 ;
        RECT 27.680 -9.370 27.950 -9.100 ;
        RECT 34.430 -9.420 34.700 -9.150 ;
        RECT 41.180 -9.370 41.450 -9.100 ;
        RECT 47.930 -9.420 48.200 -9.150 ;
        RECT 54.680 -9.370 54.950 -9.100 ;
        RECT 61.430 -9.420 61.700 -9.150 ;
        RECT 68.180 -9.370 68.450 -9.100 ;
        RECT 74.930 -9.420 75.200 -9.150 ;
        RECT 81.680 -9.370 81.950 -9.100 ;
        RECT 88.430 -9.420 88.700 -9.150 ;
        RECT 95.180 -9.370 95.450 -9.100 ;
        RECT 101.930 -9.420 102.200 -9.150 ;
        RECT 108.680 -9.370 108.950 -9.100 ;
        RECT 115.430 -9.420 115.700 -9.150 ;
        RECT 122.180 -9.370 122.450 -9.100 ;
        RECT 128.930 -9.420 129.200 -9.150 ;
        RECT 135.680 -9.370 135.950 -9.100 ;
        RECT 142.430 -9.420 142.700 -9.150 ;
        RECT 149.180 -9.370 149.450 -9.100 ;
        RECT 155.930 -9.420 156.200 -9.150 ;
        RECT 162.680 -9.370 162.950 -9.100 ;
        RECT 169.430 -9.420 169.700 -9.150 ;
        RECT 176.180 -9.370 176.450 -9.100 ;
        RECT 182.930 -9.420 183.200 -9.150 ;
        RECT 189.680 -9.370 189.950 -9.100 ;
        RECT 196.430 -9.420 196.700 -9.150 ;
        RECT 203.180 -9.370 203.450 -9.100 ;
        RECT 209.930 -9.420 210.200 -9.150 ;
        RECT 216.680 -9.370 216.950 -9.100 ;
      LAYER met2 ;
        RECT 0.590 -9.010 1.070 -9.000 ;
        RECT 108.560 -9.010 109.070 -9.000 ;
        RECT 216.560 -9.010 217.040 -9.000 ;
        RECT 0.590 -9.530 217.040 -9.010 ;
    END
  END WL14
  PIN WL15
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER li1 ;
        RECT 0.590 -10.850 1.040 -10.410 ;
        RECT 14.090 -10.850 14.540 -10.410 ;
        RECT 27.590 -10.850 28.040 -10.410 ;
        RECT 41.090 -10.850 41.540 -10.410 ;
        RECT 54.590 -10.850 55.040 -10.410 ;
        RECT 68.090 -10.850 68.540 -10.410 ;
        RECT 81.590 -10.850 82.040 -10.410 ;
        RECT 95.090 -10.850 95.540 -10.410 ;
        RECT 108.590 -10.850 109.040 -10.410 ;
        RECT 122.090 -10.850 122.540 -10.410 ;
        RECT 135.590 -10.850 136.040 -10.410 ;
        RECT 149.090 -10.850 149.540 -10.410 ;
        RECT 162.590 -10.850 163.040 -10.410 ;
        RECT 176.090 -10.850 176.540 -10.410 ;
        RECT 189.590 -10.850 190.040 -10.410 ;
        RECT 203.090 -10.850 203.540 -10.410 ;
        RECT 216.590 -10.850 217.040 -10.410 ;
        RECT 7.340 -11.770 7.790 -11.320 ;
        RECT 20.840 -11.770 21.290 -11.320 ;
        RECT 34.340 -11.770 34.790 -11.320 ;
        RECT 47.840 -11.770 48.290 -11.320 ;
        RECT 61.340 -11.770 61.790 -11.320 ;
        RECT 74.840 -11.770 75.290 -11.320 ;
        RECT 88.340 -11.770 88.790 -11.320 ;
        RECT 101.840 -11.770 102.290 -11.320 ;
        RECT 115.340 -11.770 115.790 -11.320 ;
        RECT 128.840 -11.770 129.290 -11.320 ;
        RECT 142.340 -11.770 142.790 -11.320 ;
        RECT 155.840 -11.770 156.290 -11.320 ;
        RECT 169.340 -11.770 169.790 -11.320 ;
        RECT 182.840 -11.770 183.290 -11.320 ;
        RECT 196.340 -11.770 196.790 -11.320 ;
        RECT 209.840 -11.770 210.290 -11.320 ;
      LAYER mcon ;
        RECT 0.680 -10.770 0.950 -10.500 ;
        RECT 14.180 -10.770 14.450 -10.500 ;
        RECT 27.680 -10.770 27.950 -10.500 ;
        RECT 41.180 -10.770 41.450 -10.500 ;
        RECT 54.680 -10.770 54.950 -10.500 ;
        RECT 68.180 -10.770 68.450 -10.500 ;
        RECT 81.680 -10.770 81.950 -10.500 ;
        RECT 95.180 -10.770 95.450 -10.500 ;
        RECT 108.680 -10.770 108.950 -10.500 ;
        RECT 122.180 -10.770 122.450 -10.500 ;
        RECT 135.680 -10.770 135.950 -10.500 ;
        RECT 149.180 -10.770 149.450 -10.500 ;
        RECT 162.680 -10.770 162.950 -10.500 ;
        RECT 176.180 -10.770 176.450 -10.500 ;
        RECT 189.680 -10.770 189.950 -10.500 ;
        RECT 203.180 -10.770 203.450 -10.500 ;
        RECT 216.680 -10.770 216.950 -10.500 ;
        RECT 7.440 -11.670 7.690 -11.420 ;
        RECT 20.940 -11.670 21.190 -11.420 ;
        RECT 34.440 -11.670 34.690 -11.420 ;
        RECT 47.940 -11.670 48.190 -11.420 ;
        RECT 61.440 -11.670 61.690 -11.420 ;
        RECT 74.940 -11.670 75.190 -11.420 ;
        RECT 88.440 -11.670 88.690 -11.420 ;
        RECT 101.940 -11.670 102.190 -11.420 ;
        RECT 115.440 -11.670 115.690 -11.420 ;
        RECT 128.940 -11.670 129.190 -11.420 ;
        RECT 142.440 -11.670 142.690 -11.420 ;
        RECT 155.940 -11.670 156.190 -11.420 ;
        RECT 169.440 -11.670 169.690 -11.420 ;
        RECT 182.940 -11.670 183.190 -11.420 ;
        RECT 196.440 -11.670 196.690 -11.420 ;
        RECT 209.940 -11.670 210.190 -11.420 ;
      LAYER met1 ;
        RECT 0.580 -10.850 1.040 -10.410 ;
        RECT 0.580 -10.860 1.050 -10.850 ;
        RECT 0.590 -11.330 1.050 -10.860 ;
        RECT 7.330 -11.780 7.800 -10.850 ;
        RECT 14.080 -11.330 14.550 -10.410 ;
        RECT 20.830 -11.780 21.300 -10.850 ;
        RECT 27.580 -11.330 28.050 -10.410 ;
        RECT 34.330 -11.780 34.800 -10.850 ;
        RECT 41.080 -11.330 41.550 -10.410 ;
        RECT 47.830 -11.780 48.300 -10.850 ;
        RECT 54.580 -11.330 55.050 -10.410 ;
        RECT 61.330 -11.780 61.800 -10.850 ;
        RECT 68.080 -11.330 68.550 -10.410 ;
        RECT 74.830 -11.780 75.300 -10.850 ;
        RECT 81.580 -11.330 82.050 -10.410 ;
        RECT 88.330 -11.780 88.800 -10.850 ;
        RECT 95.080 -11.330 95.550 -10.410 ;
        RECT 101.830 -11.780 102.300 -10.850 ;
        RECT 108.580 -11.330 109.050 -10.410 ;
        RECT 115.330 -11.780 115.800 -10.850 ;
        RECT 122.080 -11.330 122.550 -10.410 ;
        RECT 128.830 -11.780 129.300 -10.850 ;
        RECT 135.580 -11.330 136.050 -10.410 ;
        RECT 142.330 -11.780 142.800 -10.850 ;
        RECT 149.080 -11.330 149.550 -10.410 ;
        RECT 155.830 -11.780 156.300 -10.850 ;
        RECT 162.580 -11.330 163.050 -10.410 ;
        RECT 169.330 -11.780 169.800 -10.850 ;
        RECT 176.080 -11.330 176.550 -10.410 ;
        RECT 182.830 -11.780 183.300 -10.850 ;
        RECT 189.580 -11.330 190.050 -10.410 ;
        RECT 196.330 -11.780 196.800 -10.850 ;
        RECT 203.080 -11.330 203.550 -10.410 ;
        RECT 216.590 -10.850 217.050 -10.410 ;
        RECT 209.830 -11.780 210.300 -10.850 ;
        RECT 216.580 -10.860 217.050 -10.850 ;
        RECT 216.580 -11.330 217.040 -10.860 ;
      LAYER via ;
        RECT 0.680 -11.270 0.950 -11.000 ;
        RECT 7.430 -11.250 7.700 -10.980 ;
        RECT 14.180 -11.270 14.450 -11.000 ;
        RECT 20.930 -11.250 21.200 -10.980 ;
        RECT 27.680 -11.270 27.950 -11.000 ;
        RECT 34.430 -11.250 34.700 -10.980 ;
        RECT 41.180 -11.270 41.450 -11.000 ;
        RECT 47.930 -11.250 48.200 -10.980 ;
        RECT 54.680 -11.270 54.950 -11.000 ;
        RECT 61.430 -11.250 61.700 -10.980 ;
        RECT 68.180 -11.270 68.450 -11.000 ;
        RECT 74.930 -11.250 75.200 -10.980 ;
        RECT 81.680 -11.270 81.950 -11.000 ;
        RECT 88.430 -11.250 88.700 -10.980 ;
        RECT 95.180 -11.270 95.450 -11.000 ;
        RECT 101.930 -11.250 102.200 -10.980 ;
        RECT 108.680 -11.270 108.950 -11.000 ;
        RECT 115.430 -11.250 115.700 -10.980 ;
        RECT 122.180 -11.270 122.450 -11.000 ;
        RECT 128.930 -11.250 129.200 -10.980 ;
        RECT 135.680 -11.270 135.950 -11.000 ;
        RECT 142.430 -11.250 142.700 -10.980 ;
        RECT 149.180 -11.270 149.450 -11.000 ;
        RECT 155.930 -11.250 156.200 -10.980 ;
        RECT 162.680 -11.270 162.950 -11.000 ;
        RECT 169.430 -11.250 169.700 -10.980 ;
        RECT 176.180 -11.270 176.450 -11.000 ;
        RECT 182.930 -11.250 183.200 -10.980 ;
        RECT 189.680 -11.270 189.950 -11.000 ;
        RECT 196.430 -11.250 196.700 -10.980 ;
        RECT 203.180 -11.270 203.450 -11.000 ;
        RECT 209.930 -11.250 210.200 -10.980 ;
        RECT 216.680 -11.270 216.950 -11.000 ;
      LAYER met2 ;
        RECT 0.590 -10.860 217.040 -10.850 ;
        RECT 0.580 -11.370 217.050 -10.860 ;
    END
  END WL15
  PIN WL16
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER li1 ;
        RECT 7.340 -12.660 7.790 -12.210 ;
        RECT 20.840 -12.660 21.290 -12.210 ;
        RECT 34.340 -12.660 34.790 -12.210 ;
        RECT 47.840 -12.660 48.290 -12.210 ;
        RECT 61.340 -12.660 61.790 -12.210 ;
        RECT 74.840 -12.660 75.290 -12.210 ;
        RECT 88.340 -12.660 88.790 -12.210 ;
        RECT 101.840 -12.660 102.290 -12.210 ;
        RECT 115.340 -12.660 115.790 -12.210 ;
        RECT 128.840 -12.660 129.290 -12.210 ;
        RECT 142.340 -12.660 142.790 -12.210 ;
        RECT 155.840 -12.660 156.290 -12.210 ;
        RECT 169.340 -12.660 169.790 -12.210 ;
        RECT 182.840 -12.660 183.290 -12.210 ;
        RECT 196.340 -12.660 196.790 -12.210 ;
        RECT 209.840 -12.660 210.290 -12.210 ;
        RECT 0.590 -13.570 1.040 -13.130 ;
        RECT 14.090 -13.570 14.540 -13.130 ;
        RECT 27.590 -13.570 28.040 -13.130 ;
        RECT 41.090 -13.570 41.540 -13.130 ;
        RECT 54.590 -13.570 55.040 -13.130 ;
        RECT 68.090 -13.570 68.540 -13.130 ;
        RECT 81.590 -13.570 82.040 -13.130 ;
        RECT 95.090 -13.570 95.540 -13.130 ;
        RECT 108.590 -13.570 109.040 -13.130 ;
        RECT 122.090 -13.570 122.540 -13.130 ;
        RECT 135.590 -13.570 136.040 -13.130 ;
        RECT 149.090 -13.570 149.540 -13.130 ;
        RECT 162.590 -13.570 163.040 -13.130 ;
        RECT 176.090 -13.570 176.540 -13.130 ;
        RECT 189.590 -13.570 190.040 -13.130 ;
        RECT 203.090 -13.570 203.540 -13.130 ;
        RECT 216.590 -13.570 217.040 -13.130 ;
      LAYER mcon ;
        RECT 7.440 -12.560 7.690 -12.310 ;
        RECT 20.940 -12.560 21.190 -12.310 ;
        RECT 34.440 -12.560 34.690 -12.310 ;
        RECT 47.940 -12.560 48.190 -12.310 ;
        RECT 61.440 -12.560 61.690 -12.310 ;
        RECT 74.940 -12.560 75.190 -12.310 ;
        RECT 88.440 -12.560 88.690 -12.310 ;
        RECT 101.940 -12.560 102.190 -12.310 ;
        RECT 115.440 -12.560 115.690 -12.310 ;
        RECT 128.940 -12.560 129.190 -12.310 ;
        RECT 142.440 -12.560 142.690 -12.310 ;
        RECT 155.940 -12.560 156.190 -12.310 ;
        RECT 169.440 -12.560 169.690 -12.310 ;
        RECT 182.940 -12.560 183.190 -12.310 ;
        RECT 196.440 -12.560 196.690 -12.310 ;
        RECT 209.940 -12.560 210.190 -12.310 ;
        RECT 0.680 -13.480 0.950 -13.210 ;
        RECT 14.180 -13.480 14.450 -13.210 ;
        RECT 27.680 -13.480 27.950 -13.210 ;
        RECT 41.180 -13.480 41.450 -13.210 ;
        RECT 54.680 -13.480 54.950 -13.210 ;
        RECT 68.180 -13.480 68.450 -13.210 ;
        RECT 81.680 -13.480 81.950 -13.210 ;
        RECT 95.180 -13.480 95.450 -13.210 ;
        RECT 108.680 -13.480 108.950 -13.210 ;
        RECT 122.180 -13.480 122.450 -13.210 ;
        RECT 135.680 -13.480 135.950 -13.210 ;
        RECT 149.180 -13.480 149.450 -13.210 ;
        RECT 162.680 -13.480 162.950 -13.210 ;
        RECT 176.180 -13.480 176.450 -13.210 ;
        RECT 189.680 -13.480 189.950 -13.210 ;
        RECT 203.180 -13.480 203.450 -13.210 ;
        RECT 216.680 -13.480 216.950 -13.210 ;
      LAYER met1 ;
        RECT 0.590 -13.120 1.050 -12.650 ;
        RECT 0.580 -13.130 1.050 -13.120 ;
        RECT 7.330 -13.130 7.800 -12.200 ;
        RECT 0.580 -13.570 1.040 -13.130 ;
        RECT 14.080 -13.570 14.550 -12.650 ;
        RECT 20.830 -13.130 21.300 -12.200 ;
        RECT 27.580 -13.570 28.050 -12.650 ;
        RECT 34.330 -13.130 34.800 -12.200 ;
        RECT 41.080 -13.570 41.550 -12.650 ;
        RECT 47.830 -13.130 48.300 -12.200 ;
        RECT 54.580 -13.570 55.050 -12.650 ;
        RECT 61.330 -13.130 61.800 -12.200 ;
        RECT 68.080 -13.570 68.550 -12.650 ;
        RECT 74.830 -13.130 75.300 -12.200 ;
        RECT 81.580 -13.570 82.050 -12.650 ;
        RECT 88.330 -13.130 88.800 -12.200 ;
        RECT 95.080 -13.570 95.550 -12.650 ;
        RECT 101.830 -13.130 102.300 -12.200 ;
        RECT 108.580 -13.570 109.050 -12.650 ;
        RECT 115.330 -13.130 115.800 -12.200 ;
        RECT 122.080 -13.570 122.550 -12.650 ;
        RECT 128.830 -13.130 129.300 -12.200 ;
        RECT 135.580 -13.570 136.050 -12.650 ;
        RECT 142.330 -13.130 142.800 -12.200 ;
        RECT 149.080 -13.570 149.550 -12.650 ;
        RECT 155.830 -13.130 156.300 -12.200 ;
        RECT 162.580 -13.570 163.050 -12.650 ;
        RECT 169.330 -13.130 169.800 -12.200 ;
        RECT 176.080 -13.570 176.550 -12.650 ;
        RECT 182.830 -13.130 183.300 -12.200 ;
        RECT 189.580 -13.570 190.050 -12.650 ;
        RECT 196.330 -13.130 196.800 -12.200 ;
        RECT 203.080 -13.570 203.550 -12.650 ;
        RECT 209.830 -13.130 210.300 -12.200 ;
        RECT 216.580 -13.120 217.040 -12.650 ;
        RECT 216.580 -13.130 217.050 -13.120 ;
        RECT 216.590 -13.570 217.050 -13.130 ;
      LAYER via ;
        RECT 0.680 -12.980 0.950 -12.710 ;
        RECT 7.430 -13.000 7.700 -12.730 ;
        RECT 14.180 -12.980 14.450 -12.710 ;
        RECT 20.930 -13.000 21.200 -12.730 ;
        RECT 27.680 -12.980 27.950 -12.710 ;
        RECT 34.430 -13.000 34.700 -12.730 ;
        RECT 41.180 -12.980 41.450 -12.710 ;
        RECT 47.930 -13.000 48.200 -12.730 ;
        RECT 54.680 -12.980 54.950 -12.710 ;
        RECT 61.430 -13.000 61.700 -12.730 ;
        RECT 68.180 -12.980 68.450 -12.710 ;
        RECT 74.930 -13.000 75.200 -12.730 ;
        RECT 81.680 -12.980 81.950 -12.710 ;
        RECT 88.430 -13.000 88.700 -12.730 ;
        RECT 95.180 -12.980 95.450 -12.710 ;
        RECT 101.930 -13.000 102.200 -12.730 ;
        RECT 108.680 -12.980 108.950 -12.710 ;
        RECT 115.430 -13.000 115.700 -12.730 ;
        RECT 122.180 -12.980 122.450 -12.710 ;
        RECT 128.930 -13.000 129.200 -12.730 ;
        RECT 135.680 -12.980 135.950 -12.710 ;
        RECT 142.430 -13.000 142.700 -12.730 ;
        RECT 149.180 -12.980 149.450 -12.710 ;
        RECT 155.930 -13.000 156.200 -12.730 ;
        RECT 162.680 -12.980 162.950 -12.710 ;
        RECT 169.430 -13.000 169.700 -12.730 ;
        RECT 176.180 -12.980 176.450 -12.710 ;
        RECT 182.930 -13.000 183.200 -12.730 ;
        RECT 189.680 -12.980 189.950 -12.710 ;
        RECT 196.430 -13.000 196.700 -12.730 ;
        RECT 203.180 -12.980 203.450 -12.710 ;
        RECT 209.930 -13.000 210.200 -12.730 ;
        RECT 216.680 -12.980 216.950 -12.710 ;
      LAYER met2 ;
        RECT 0.580 -13.120 217.050 -12.610 ;
        RECT 0.590 -13.130 217.040 -13.120 ;
    END
  END WL16
  PIN WL17
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER li1 ;
        RECT 0.590 -14.460 1.040 -14.020 ;
        RECT 14.090 -14.460 14.540 -14.020 ;
        RECT 27.590 -14.460 28.040 -14.020 ;
        RECT 41.090 -14.460 41.540 -14.020 ;
        RECT 54.590 -14.460 55.040 -14.020 ;
        RECT 68.090 -14.460 68.540 -14.020 ;
        RECT 81.590 -14.460 82.040 -14.020 ;
        RECT 95.090 -14.460 95.540 -14.020 ;
        RECT 108.590 -14.460 109.040 -14.020 ;
        RECT 122.090 -14.460 122.540 -14.020 ;
        RECT 135.590 -14.460 136.040 -14.020 ;
        RECT 149.090 -14.460 149.540 -14.020 ;
        RECT 162.590 -14.460 163.040 -14.020 ;
        RECT 176.090 -14.460 176.540 -14.020 ;
        RECT 189.590 -14.460 190.040 -14.020 ;
        RECT 203.090 -14.460 203.540 -14.020 ;
        RECT 216.590 -14.460 217.040 -14.020 ;
        RECT 7.340 -15.380 7.790 -14.930 ;
        RECT 20.840 -15.380 21.290 -14.930 ;
        RECT 34.340 -15.380 34.790 -14.930 ;
        RECT 47.840 -15.380 48.290 -14.930 ;
        RECT 61.340 -15.380 61.790 -14.930 ;
        RECT 74.840 -15.380 75.290 -14.930 ;
        RECT 88.340 -15.380 88.790 -14.930 ;
        RECT 101.840 -15.380 102.290 -14.930 ;
        RECT 115.340 -15.380 115.790 -14.930 ;
        RECT 128.840 -15.380 129.290 -14.930 ;
        RECT 142.340 -15.380 142.790 -14.930 ;
        RECT 155.840 -15.380 156.290 -14.930 ;
        RECT 169.340 -15.380 169.790 -14.930 ;
        RECT 182.840 -15.380 183.290 -14.930 ;
        RECT 196.340 -15.380 196.790 -14.930 ;
        RECT 209.840 -15.380 210.290 -14.930 ;
      LAYER mcon ;
        RECT 0.680 -14.380 0.950 -14.110 ;
        RECT 14.180 -14.380 14.450 -14.110 ;
        RECT 27.680 -14.380 27.950 -14.110 ;
        RECT 41.180 -14.380 41.450 -14.110 ;
        RECT 54.680 -14.380 54.950 -14.110 ;
        RECT 68.180 -14.380 68.450 -14.110 ;
        RECT 81.680 -14.380 81.950 -14.110 ;
        RECT 95.180 -14.380 95.450 -14.110 ;
        RECT 108.680 -14.380 108.950 -14.110 ;
        RECT 122.180 -14.380 122.450 -14.110 ;
        RECT 135.680 -14.380 135.950 -14.110 ;
        RECT 149.180 -14.380 149.450 -14.110 ;
        RECT 162.680 -14.380 162.950 -14.110 ;
        RECT 176.180 -14.380 176.450 -14.110 ;
        RECT 189.680 -14.380 189.950 -14.110 ;
        RECT 203.180 -14.380 203.450 -14.110 ;
        RECT 216.680 -14.380 216.950 -14.110 ;
        RECT 7.440 -15.280 7.690 -15.030 ;
        RECT 20.940 -15.280 21.190 -15.030 ;
        RECT 34.440 -15.280 34.690 -15.030 ;
        RECT 47.940 -15.280 48.190 -15.030 ;
        RECT 61.440 -15.280 61.690 -15.030 ;
        RECT 74.940 -15.280 75.190 -15.030 ;
        RECT 88.440 -15.280 88.690 -15.030 ;
        RECT 101.940 -15.280 102.190 -15.030 ;
        RECT 115.440 -15.280 115.690 -15.030 ;
        RECT 128.940 -15.280 129.190 -15.030 ;
        RECT 142.440 -15.280 142.690 -15.030 ;
        RECT 155.940 -15.280 156.190 -15.030 ;
        RECT 169.440 -15.280 169.690 -15.030 ;
        RECT 182.940 -15.280 183.190 -15.030 ;
        RECT 196.440 -15.280 196.690 -15.030 ;
        RECT 209.940 -15.280 210.190 -15.030 ;
      LAYER met1 ;
        RECT 0.580 -14.460 1.040 -14.020 ;
        RECT 0.580 -14.470 1.050 -14.460 ;
        RECT 0.590 -14.940 1.050 -14.470 ;
        RECT 7.330 -15.390 7.800 -14.460 ;
        RECT 14.080 -14.940 14.550 -14.020 ;
        RECT 20.830 -15.390 21.300 -14.460 ;
        RECT 27.580 -14.940 28.050 -14.020 ;
        RECT 34.330 -15.390 34.800 -14.460 ;
        RECT 41.080 -14.940 41.550 -14.020 ;
        RECT 47.830 -15.390 48.300 -14.460 ;
        RECT 54.580 -14.940 55.050 -14.020 ;
        RECT 61.330 -15.390 61.800 -14.460 ;
        RECT 68.080 -14.940 68.550 -14.020 ;
        RECT 74.830 -15.390 75.300 -14.460 ;
        RECT 81.580 -14.940 82.050 -14.020 ;
        RECT 88.330 -15.390 88.800 -14.460 ;
        RECT 95.080 -14.940 95.550 -14.020 ;
        RECT 101.830 -15.390 102.300 -14.460 ;
        RECT 108.580 -14.940 109.050 -14.020 ;
        RECT 115.330 -15.390 115.800 -14.460 ;
        RECT 122.080 -14.940 122.550 -14.020 ;
        RECT 128.830 -15.390 129.300 -14.460 ;
        RECT 135.580 -14.940 136.050 -14.020 ;
        RECT 142.330 -15.390 142.800 -14.460 ;
        RECT 149.080 -14.940 149.550 -14.020 ;
        RECT 155.830 -15.390 156.300 -14.460 ;
        RECT 162.580 -14.940 163.050 -14.020 ;
        RECT 169.330 -15.390 169.800 -14.460 ;
        RECT 176.080 -14.940 176.550 -14.020 ;
        RECT 182.830 -15.390 183.300 -14.460 ;
        RECT 189.580 -14.940 190.050 -14.020 ;
        RECT 196.330 -15.390 196.800 -14.460 ;
        RECT 203.080 -14.940 203.550 -14.020 ;
        RECT 216.590 -14.460 217.050 -14.020 ;
        RECT 209.830 -15.390 210.300 -14.460 ;
        RECT 216.580 -14.470 217.050 -14.460 ;
        RECT 216.580 -14.940 217.040 -14.470 ;
      LAYER via ;
        RECT 0.680 -14.880 0.950 -14.610 ;
        RECT 7.430 -14.830 7.700 -14.560 ;
        RECT 14.180 -14.880 14.450 -14.610 ;
        RECT 20.930 -14.830 21.200 -14.560 ;
        RECT 27.680 -14.880 27.950 -14.610 ;
        RECT 34.430 -14.830 34.700 -14.560 ;
        RECT 41.180 -14.880 41.450 -14.610 ;
        RECT 47.930 -14.830 48.200 -14.560 ;
        RECT 54.680 -14.880 54.950 -14.610 ;
        RECT 61.430 -14.830 61.700 -14.560 ;
        RECT 68.180 -14.880 68.450 -14.610 ;
        RECT 74.930 -14.830 75.200 -14.560 ;
        RECT 81.680 -14.880 81.950 -14.610 ;
        RECT 88.430 -14.830 88.700 -14.560 ;
        RECT 95.180 -14.880 95.450 -14.610 ;
        RECT 101.930 -14.830 102.200 -14.560 ;
        RECT 108.680 -14.880 108.950 -14.610 ;
        RECT 115.430 -14.830 115.700 -14.560 ;
        RECT 122.180 -14.880 122.450 -14.610 ;
        RECT 128.930 -14.830 129.200 -14.560 ;
        RECT 135.680 -14.880 135.950 -14.610 ;
        RECT 142.430 -14.830 142.700 -14.560 ;
        RECT 149.180 -14.880 149.450 -14.610 ;
        RECT 155.930 -14.830 156.200 -14.560 ;
        RECT 162.680 -14.880 162.950 -14.610 ;
        RECT 169.430 -14.830 169.700 -14.560 ;
        RECT 176.180 -14.880 176.450 -14.610 ;
        RECT 182.930 -14.830 183.200 -14.560 ;
        RECT 189.680 -14.880 189.950 -14.610 ;
        RECT 196.430 -14.830 196.700 -14.560 ;
        RECT 203.180 -14.880 203.450 -14.610 ;
        RECT 209.930 -14.830 210.200 -14.560 ;
        RECT 216.680 -14.880 216.950 -14.610 ;
      LAYER met2 ;
        RECT 0.590 -14.970 217.040 -14.450 ;
        RECT 0.590 -14.980 1.070 -14.970 ;
        RECT 108.560 -14.980 109.070 -14.970 ;
        RECT 216.560 -14.980 217.040 -14.970 ;
    END
  END WL17
  PIN WL18
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER li1 ;
        RECT 7.340 -16.270 7.790 -15.820 ;
        RECT 20.840 -16.270 21.290 -15.820 ;
        RECT 34.340 -16.270 34.790 -15.820 ;
        RECT 47.840 -16.270 48.290 -15.820 ;
        RECT 61.340 -16.270 61.790 -15.820 ;
        RECT 74.840 -16.270 75.290 -15.820 ;
        RECT 88.340 -16.270 88.790 -15.820 ;
        RECT 101.840 -16.270 102.290 -15.820 ;
        RECT 115.340 -16.270 115.790 -15.820 ;
        RECT 128.840 -16.270 129.290 -15.820 ;
        RECT 142.340 -16.270 142.790 -15.820 ;
        RECT 155.840 -16.270 156.290 -15.820 ;
        RECT 169.340 -16.270 169.790 -15.820 ;
        RECT 182.840 -16.270 183.290 -15.820 ;
        RECT 196.340 -16.270 196.790 -15.820 ;
        RECT 209.840 -16.270 210.290 -15.820 ;
        RECT 0.590 -17.180 1.040 -16.740 ;
        RECT 14.090 -17.180 14.540 -16.740 ;
        RECT 27.590 -17.180 28.040 -16.740 ;
        RECT 41.090 -17.180 41.540 -16.740 ;
        RECT 54.590 -17.180 55.040 -16.740 ;
        RECT 68.090 -17.180 68.540 -16.740 ;
        RECT 81.590 -17.180 82.040 -16.740 ;
        RECT 95.090 -17.180 95.540 -16.740 ;
        RECT 108.590 -17.180 109.040 -16.740 ;
        RECT 122.090 -17.180 122.540 -16.740 ;
        RECT 135.590 -17.180 136.040 -16.740 ;
        RECT 149.090 -17.180 149.540 -16.740 ;
        RECT 162.590 -17.180 163.040 -16.740 ;
        RECT 176.090 -17.180 176.540 -16.740 ;
        RECT 189.590 -17.180 190.040 -16.740 ;
        RECT 203.090 -17.180 203.540 -16.740 ;
        RECT 216.590 -17.180 217.040 -16.740 ;
      LAYER mcon ;
        RECT 7.440 -16.170 7.690 -15.920 ;
        RECT 20.940 -16.170 21.190 -15.920 ;
        RECT 34.440 -16.170 34.690 -15.920 ;
        RECT 47.940 -16.170 48.190 -15.920 ;
        RECT 61.440 -16.170 61.690 -15.920 ;
        RECT 74.940 -16.170 75.190 -15.920 ;
        RECT 88.440 -16.170 88.690 -15.920 ;
        RECT 101.940 -16.170 102.190 -15.920 ;
        RECT 115.440 -16.170 115.690 -15.920 ;
        RECT 128.940 -16.170 129.190 -15.920 ;
        RECT 142.440 -16.170 142.690 -15.920 ;
        RECT 155.940 -16.170 156.190 -15.920 ;
        RECT 169.440 -16.170 169.690 -15.920 ;
        RECT 182.940 -16.170 183.190 -15.920 ;
        RECT 196.440 -16.170 196.690 -15.920 ;
        RECT 209.940 -16.170 210.190 -15.920 ;
        RECT 0.680 -17.090 0.950 -16.820 ;
        RECT 14.180 -17.090 14.450 -16.820 ;
        RECT 27.680 -17.090 27.950 -16.820 ;
        RECT 41.180 -17.090 41.450 -16.820 ;
        RECT 54.680 -17.090 54.950 -16.820 ;
        RECT 68.180 -17.090 68.450 -16.820 ;
        RECT 81.680 -17.090 81.950 -16.820 ;
        RECT 95.180 -17.090 95.450 -16.820 ;
        RECT 108.680 -17.090 108.950 -16.820 ;
        RECT 122.180 -17.090 122.450 -16.820 ;
        RECT 135.680 -17.090 135.950 -16.820 ;
        RECT 149.180 -17.090 149.450 -16.820 ;
        RECT 162.680 -17.090 162.950 -16.820 ;
        RECT 176.180 -17.090 176.450 -16.820 ;
        RECT 189.680 -17.090 189.950 -16.820 ;
        RECT 203.180 -17.090 203.450 -16.820 ;
        RECT 216.680 -17.090 216.950 -16.820 ;
      LAYER met1 ;
        RECT 0.590 -16.730 1.050 -16.260 ;
        RECT 0.580 -16.740 1.050 -16.730 ;
        RECT 7.330 -16.740 7.800 -15.810 ;
        RECT 0.580 -17.180 1.040 -16.740 ;
        RECT 14.080 -17.180 14.550 -16.260 ;
        RECT 20.830 -16.740 21.300 -15.810 ;
        RECT 27.580 -17.180 28.050 -16.260 ;
        RECT 34.330 -16.740 34.800 -15.810 ;
        RECT 41.080 -17.180 41.550 -16.260 ;
        RECT 47.830 -16.740 48.300 -15.810 ;
        RECT 54.580 -17.180 55.050 -16.260 ;
        RECT 61.330 -16.740 61.800 -15.810 ;
        RECT 68.080 -17.180 68.550 -16.260 ;
        RECT 74.830 -16.740 75.300 -15.810 ;
        RECT 81.580 -17.180 82.050 -16.260 ;
        RECT 88.330 -16.740 88.800 -15.810 ;
        RECT 95.080 -17.180 95.550 -16.260 ;
        RECT 101.830 -16.740 102.300 -15.810 ;
        RECT 108.580 -17.180 109.050 -16.260 ;
        RECT 115.330 -16.740 115.800 -15.810 ;
        RECT 122.080 -17.180 122.550 -16.260 ;
        RECT 128.830 -16.740 129.300 -15.810 ;
        RECT 135.580 -17.180 136.050 -16.260 ;
        RECT 142.330 -16.740 142.800 -15.810 ;
        RECT 149.080 -17.180 149.550 -16.260 ;
        RECT 155.830 -16.740 156.300 -15.810 ;
        RECT 162.580 -17.180 163.050 -16.260 ;
        RECT 169.330 -16.740 169.800 -15.810 ;
        RECT 176.080 -17.180 176.550 -16.260 ;
        RECT 182.830 -16.740 183.300 -15.810 ;
        RECT 189.580 -17.180 190.050 -16.260 ;
        RECT 196.330 -16.740 196.800 -15.810 ;
        RECT 203.080 -17.180 203.550 -16.260 ;
        RECT 209.830 -16.740 210.300 -15.810 ;
        RECT 216.580 -16.730 217.040 -16.260 ;
        RECT 216.580 -16.740 217.050 -16.730 ;
        RECT 216.590 -17.180 217.050 -16.740 ;
      LAYER via ;
        RECT 0.680 -16.590 0.950 -16.320 ;
        RECT 7.430 -16.610 7.700 -16.340 ;
        RECT 14.180 -16.590 14.450 -16.320 ;
        RECT 20.930 -16.640 21.200 -16.370 ;
        RECT 27.680 -16.590 27.950 -16.320 ;
        RECT 34.430 -16.640 34.700 -16.370 ;
        RECT 41.180 -16.590 41.450 -16.320 ;
        RECT 47.930 -16.610 48.200 -16.340 ;
        RECT 54.680 -16.590 54.950 -16.320 ;
        RECT 61.430 -16.610 61.700 -16.340 ;
        RECT 68.180 -16.590 68.450 -16.320 ;
        RECT 74.930 -16.640 75.200 -16.370 ;
        RECT 81.680 -16.590 81.950 -16.320 ;
        RECT 88.430 -16.640 88.700 -16.370 ;
        RECT 95.180 -16.590 95.450 -16.320 ;
        RECT 101.930 -16.610 102.200 -16.340 ;
        RECT 108.680 -16.590 108.950 -16.320 ;
        RECT 115.430 -16.610 115.700 -16.340 ;
        RECT 122.180 -16.590 122.450 -16.320 ;
        RECT 128.930 -16.640 129.200 -16.370 ;
        RECT 135.680 -16.590 135.950 -16.320 ;
        RECT 142.430 -16.640 142.700 -16.370 ;
        RECT 149.180 -16.590 149.450 -16.320 ;
        RECT 155.930 -16.610 156.200 -16.340 ;
        RECT 162.680 -16.590 162.950 -16.320 ;
        RECT 169.430 -16.610 169.700 -16.340 ;
        RECT 176.180 -16.590 176.450 -16.320 ;
        RECT 182.930 -16.640 183.200 -16.370 ;
        RECT 189.680 -16.590 189.950 -16.320 ;
        RECT 196.430 -16.640 196.700 -16.370 ;
        RECT 203.180 -16.590 203.450 -16.320 ;
        RECT 209.930 -16.610 210.200 -16.340 ;
        RECT 216.680 -16.590 216.950 -16.320 ;
      LAYER met2 ;
        RECT 0.590 -16.220 1.070 -16.210 ;
        RECT 108.560 -16.220 109.070 -16.210 ;
        RECT 216.560 -16.220 217.040 -16.210 ;
        RECT 0.590 -16.230 14.590 -16.220 ;
        RECT 41.040 -16.230 68.590 -16.220 ;
        RECT 95.040 -16.230 122.590 -16.220 ;
        RECT 149.040 -16.230 176.590 -16.220 ;
        RECT 203.040 -16.230 217.040 -16.220 ;
        RECT 0.590 -16.250 217.040 -16.230 ;
        RECT 0.580 -16.730 217.050 -16.250 ;
        RECT 0.590 -16.740 217.040 -16.730 ;
        RECT 14.040 -16.750 41.590 -16.740 ;
        RECT 68.040 -16.750 95.590 -16.740 ;
        RECT 122.040 -16.750 149.590 -16.740 ;
        RECT 176.040 -16.750 203.590 -16.740 ;
    END
  END WL18
  PIN WL19
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER li1 ;
        RECT 0.590 -18.070 1.040 -17.630 ;
        RECT 14.090 -18.070 14.540 -17.630 ;
        RECT 27.590 -18.070 28.040 -17.630 ;
        RECT 41.090 -18.070 41.540 -17.630 ;
        RECT 54.590 -18.070 55.040 -17.630 ;
        RECT 68.090 -18.070 68.540 -17.630 ;
        RECT 81.590 -18.070 82.040 -17.630 ;
        RECT 95.090 -18.070 95.540 -17.630 ;
        RECT 108.590 -18.070 109.040 -17.630 ;
        RECT 122.090 -18.070 122.540 -17.630 ;
        RECT 135.590 -18.070 136.040 -17.630 ;
        RECT 149.090 -18.070 149.540 -17.630 ;
        RECT 162.590 -18.070 163.040 -17.630 ;
        RECT 176.090 -18.070 176.540 -17.630 ;
        RECT 189.590 -18.070 190.040 -17.630 ;
        RECT 203.090 -18.070 203.540 -17.630 ;
        RECT 216.590 -18.070 217.040 -17.630 ;
        RECT 7.340 -18.990 7.790 -18.540 ;
        RECT 20.840 -18.990 21.290 -18.540 ;
        RECT 34.340 -18.990 34.790 -18.540 ;
        RECT 47.840 -18.990 48.290 -18.540 ;
        RECT 61.340 -18.990 61.790 -18.540 ;
        RECT 74.840 -18.990 75.290 -18.540 ;
        RECT 88.340 -18.990 88.790 -18.540 ;
        RECT 101.840 -18.990 102.290 -18.540 ;
        RECT 115.340 -18.990 115.790 -18.540 ;
        RECT 128.840 -18.990 129.290 -18.540 ;
        RECT 142.340 -18.990 142.790 -18.540 ;
        RECT 155.840 -18.990 156.290 -18.540 ;
        RECT 169.340 -18.990 169.790 -18.540 ;
        RECT 182.840 -18.990 183.290 -18.540 ;
        RECT 196.340 -18.990 196.790 -18.540 ;
        RECT 209.840 -18.990 210.290 -18.540 ;
      LAYER mcon ;
        RECT 0.680 -17.990 0.950 -17.720 ;
        RECT 14.180 -17.990 14.450 -17.720 ;
        RECT 27.680 -17.990 27.950 -17.720 ;
        RECT 41.180 -17.990 41.450 -17.720 ;
        RECT 54.680 -17.990 54.950 -17.720 ;
        RECT 68.180 -17.990 68.450 -17.720 ;
        RECT 81.680 -17.990 81.950 -17.720 ;
        RECT 95.180 -17.990 95.450 -17.720 ;
        RECT 108.680 -17.990 108.950 -17.720 ;
        RECT 122.180 -17.990 122.450 -17.720 ;
        RECT 135.680 -17.990 135.950 -17.720 ;
        RECT 149.180 -17.990 149.450 -17.720 ;
        RECT 162.680 -17.990 162.950 -17.720 ;
        RECT 176.180 -17.990 176.450 -17.720 ;
        RECT 189.680 -17.990 189.950 -17.720 ;
        RECT 203.180 -17.990 203.450 -17.720 ;
        RECT 216.680 -17.990 216.950 -17.720 ;
        RECT 7.440 -18.890 7.690 -18.640 ;
        RECT 20.940 -18.890 21.190 -18.640 ;
        RECT 34.440 -18.890 34.690 -18.640 ;
        RECT 47.940 -18.890 48.190 -18.640 ;
        RECT 61.440 -18.890 61.690 -18.640 ;
        RECT 74.940 -18.890 75.190 -18.640 ;
        RECT 88.440 -18.890 88.690 -18.640 ;
        RECT 101.940 -18.890 102.190 -18.640 ;
        RECT 115.440 -18.890 115.690 -18.640 ;
        RECT 128.940 -18.890 129.190 -18.640 ;
        RECT 142.440 -18.890 142.690 -18.640 ;
        RECT 155.940 -18.890 156.190 -18.640 ;
        RECT 169.440 -18.890 169.690 -18.640 ;
        RECT 182.940 -18.890 183.190 -18.640 ;
        RECT 196.440 -18.890 196.690 -18.640 ;
        RECT 209.940 -18.890 210.190 -18.640 ;
      LAYER met1 ;
        RECT 0.580 -18.070 1.040 -17.630 ;
        RECT 0.580 -18.080 1.050 -18.070 ;
        RECT 0.590 -18.550 1.050 -18.080 ;
        RECT 7.330 -19.000 7.800 -18.070 ;
        RECT 14.080 -18.550 14.550 -17.630 ;
        RECT 20.830 -19.000 21.300 -18.070 ;
        RECT 27.580 -18.550 28.050 -17.630 ;
        RECT 34.330 -19.000 34.800 -18.070 ;
        RECT 41.080 -18.550 41.550 -17.630 ;
        RECT 47.830 -19.000 48.300 -18.070 ;
        RECT 54.580 -18.550 55.050 -17.630 ;
        RECT 61.330 -19.000 61.800 -18.070 ;
        RECT 68.080 -18.550 68.550 -17.630 ;
        RECT 74.830 -19.000 75.300 -18.070 ;
        RECT 81.580 -18.550 82.050 -17.630 ;
        RECT 88.330 -19.000 88.800 -18.070 ;
        RECT 95.080 -18.550 95.550 -17.630 ;
        RECT 101.830 -19.000 102.300 -18.070 ;
        RECT 108.580 -18.550 109.050 -17.630 ;
        RECT 115.330 -19.000 115.800 -18.070 ;
        RECT 122.080 -18.550 122.550 -17.630 ;
        RECT 128.830 -19.000 129.300 -18.070 ;
        RECT 135.580 -18.550 136.050 -17.630 ;
        RECT 142.330 -19.000 142.800 -18.070 ;
        RECT 149.080 -18.550 149.550 -17.630 ;
        RECT 155.830 -19.000 156.300 -18.070 ;
        RECT 162.580 -18.550 163.050 -17.630 ;
        RECT 169.330 -19.000 169.800 -18.070 ;
        RECT 176.080 -18.550 176.550 -17.630 ;
        RECT 182.830 -19.000 183.300 -18.070 ;
        RECT 189.580 -18.550 190.050 -17.630 ;
        RECT 196.330 -19.000 196.800 -18.070 ;
        RECT 203.080 -18.550 203.550 -17.630 ;
        RECT 216.590 -18.070 217.050 -17.630 ;
        RECT 209.830 -19.000 210.300 -18.070 ;
        RECT 216.580 -18.080 217.050 -18.070 ;
        RECT 216.580 -18.550 217.040 -18.080 ;
      LAYER via ;
        RECT 0.680 -18.490 0.950 -18.220 ;
        RECT 7.430 -18.440 7.700 -18.170 ;
        RECT 14.180 -18.490 14.450 -18.220 ;
        RECT 20.930 -18.470 21.200 -18.200 ;
        RECT 27.680 -18.490 27.950 -18.220 ;
        RECT 34.430 -18.470 34.700 -18.200 ;
        RECT 41.180 -18.490 41.450 -18.220 ;
        RECT 47.930 -18.440 48.200 -18.170 ;
        RECT 54.680 -18.490 54.950 -18.220 ;
        RECT 61.430 -18.440 61.700 -18.170 ;
        RECT 68.180 -18.490 68.450 -18.220 ;
        RECT 74.930 -18.470 75.200 -18.200 ;
        RECT 81.680 -18.490 81.950 -18.220 ;
        RECT 88.430 -18.470 88.700 -18.200 ;
        RECT 95.180 -18.490 95.450 -18.220 ;
        RECT 101.930 -18.440 102.200 -18.170 ;
        RECT 108.680 -18.490 108.950 -18.220 ;
        RECT 115.430 -18.440 115.700 -18.170 ;
        RECT 122.180 -18.490 122.450 -18.220 ;
        RECT 128.930 -18.470 129.200 -18.200 ;
        RECT 135.680 -18.490 135.950 -18.220 ;
        RECT 142.430 -18.470 142.700 -18.200 ;
        RECT 149.180 -18.490 149.450 -18.220 ;
        RECT 155.930 -18.440 156.200 -18.170 ;
        RECT 162.680 -18.490 162.950 -18.220 ;
        RECT 169.430 -18.440 169.700 -18.170 ;
        RECT 176.180 -18.490 176.450 -18.220 ;
        RECT 182.930 -18.470 183.200 -18.200 ;
        RECT 189.680 -18.490 189.950 -18.220 ;
        RECT 196.430 -18.470 196.700 -18.200 ;
        RECT 203.180 -18.490 203.450 -18.220 ;
        RECT 209.930 -18.440 210.200 -18.170 ;
        RECT 216.680 -18.490 216.950 -18.220 ;
      LAYER met2 ;
        RECT 0.590 -18.070 14.590 -18.060 ;
        RECT 41.040 -18.070 68.590 -18.060 ;
        RECT 95.040 -18.070 122.590 -18.060 ;
        RECT 149.040 -18.070 176.590 -18.060 ;
        RECT 203.040 -18.070 217.040 -18.060 ;
        RECT 0.590 -18.090 217.040 -18.070 ;
        RECT 0.580 -18.570 217.050 -18.090 ;
        RECT 0.590 -18.580 217.040 -18.570 ;
        RECT 14.040 -18.590 41.590 -18.580 ;
        RECT 68.040 -18.590 95.590 -18.580 ;
        RECT 122.040 -18.590 149.590 -18.580 ;
        RECT 176.040 -18.590 203.590 -18.580 ;
    END
  END WL19
  PIN WL20
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER li1 ;
        RECT 7.340 -19.880 7.790 -19.430 ;
        RECT 20.840 -19.880 21.290 -19.430 ;
        RECT 34.340 -19.880 34.790 -19.430 ;
        RECT 47.840 -19.880 48.290 -19.430 ;
        RECT 61.340 -19.880 61.790 -19.430 ;
        RECT 74.840 -19.880 75.290 -19.430 ;
        RECT 88.340 -19.880 88.790 -19.430 ;
        RECT 101.840 -19.880 102.290 -19.430 ;
        RECT 115.340 -19.880 115.790 -19.430 ;
        RECT 128.840 -19.880 129.290 -19.430 ;
        RECT 142.340 -19.880 142.790 -19.430 ;
        RECT 155.840 -19.880 156.290 -19.430 ;
        RECT 169.340 -19.880 169.790 -19.430 ;
        RECT 182.840 -19.880 183.290 -19.430 ;
        RECT 196.340 -19.880 196.790 -19.430 ;
        RECT 209.840 -19.880 210.290 -19.430 ;
        RECT 0.590 -20.790 1.040 -20.350 ;
        RECT 14.090 -20.790 14.540 -20.350 ;
        RECT 27.590 -20.790 28.040 -20.350 ;
        RECT 41.090 -20.790 41.540 -20.350 ;
        RECT 54.590 -20.790 55.040 -20.350 ;
        RECT 68.090 -20.790 68.540 -20.350 ;
        RECT 81.590 -20.790 82.040 -20.350 ;
        RECT 95.090 -20.790 95.540 -20.350 ;
        RECT 108.590 -20.790 109.040 -20.350 ;
        RECT 122.090 -20.790 122.540 -20.350 ;
        RECT 135.590 -20.790 136.040 -20.350 ;
        RECT 149.090 -20.790 149.540 -20.350 ;
        RECT 162.590 -20.790 163.040 -20.350 ;
        RECT 176.090 -20.790 176.540 -20.350 ;
        RECT 189.590 -20.790 190.040 -20.350 ;
        RECT 203.090 -20.790 203.540 -20.350 ;
        RECT 216.590 -20.790 217.040 -20.350 ;
      LAYER mcon ;
        RECT 7.440 -19.780 7.690 -19.530 ;
        RECT 20.940 -19.780 21.190 -19.530 ;
        RECT 34.440 -19.780 34.690 -19.530 ;
        RECT 47.940 -19.780 48.190 -19.530 ;
        RECT 61.440 -19.780 61.690 -19.530 ;
        RECT 74.940 -19.780 75.190 -19.530 ;
        RECT 88.440 -19.780 88.690 -19.530 ;
        RECT 101.940 -19.780 102.190 -19.530 ;
        RECT 115.440 -19.780 115.690 -19.530 ;
        RECT 128.940 -19.780 129.190 -19.530 ;
        RECT 142.440 -19.780 142.690 -19.530 ;
        RECT 155.940 -19.780 156.190 -19.530 ;
        RECT 169.440 -19.780 169.690 -19.530 ;
        RECT 182.940 -19.780 183.190 -19.530 ;
        RECT 196.440 -19.780 196.690 -19.530 ;
        RECT 209.940 -19.780 210.190 -19.530 ;
        RECT 0.680 -20.700 0.950 -20.430 ;
        RECT 14.180 -20.700 14.450 -20.430 ;
        RECT 27.680 -20.700 27.950 -20.430 ;
        RECT 41.180 -20.700 41.450 -20.430 ;
        RECT 54.680 -20.700 54.950 -20.430 ;
        RECT 68.180 -20.700 68.450 -20.430 ;
        RECT 81.680 -20.700 81.950 -20.430 ;
        RECT 95.180 -20.700 95.450 -20.430 ;
        RECT 108.680 -20.700 108.950 -20.430 ;
        RECT 122.180 -20.700 122.450 -20.430 ;
        RECT 135.680 -20.700 135.950 -20.430 ;
        RECT 149.180 -20.700 149.450 -20.430 ;
        RECT 162.680 -20.700 162.950 -20.430 ;
        RECT 176.180 -20.700 176.450 -20.430 ;
        RECT 189.680 -20.700 189.950 -20.430 ;
        RECT 203.180 -20.700 203.450 -20.430 ;
        RECT 216.680 -20.700 216.950 -20.430 ;
      LAYER met1 ;
        RECT 0.590 -20.340 1.050 -19.870 ;
        RECT 0.580 -20.350 1.050 -20.340 ;
        RECT 7.330 -20.350 7.800 -19.420 ;
        RECT 0.580 -20.790 1.040 -20.350 ;
        RECT 14.080 -20.790 14.550 -19.870 ;
        RECT 20.830 -20.350 21.300 -19.420 ;
        RECT 27.580 -20.790 28.050 -19.870 ;
        RECT 34.330 -20.350 34.800 -19.420 ;
        RECT 41.080 -20.790 41.550 -19.870 ;
        RECT 47.830 -20.350 48.300 -19.420 ;
        RECT 54.580 -20.790 55.050 -19.870 ;
        RECT 61.330 -20.350 61.800 -19.420 ;
        RECT 68.080 -20.790 68.550 -19.870 ;
        RECT 74.830 -20.350 75.300 -19.420 ;
        RECT 81.580 -20.790 82.050 -19.870 ;
        RECT 88.330 -20.350 88.800 -19.420 ;
        RECT 95.080 -20.790 95.550 -19.870 ;
        RECT 101.830 -20.350 102.300 -19.420 ;
        RECT 108.580 -20.790 109.050 -19.870 ;
        RECT 115.330 -20.350 115.800 -19.420 ;
        RECT 122.080 -20.790 122.550 -19.870 ;
        RECT 128.830 -20.350 129.300 -19.420 ;
        RECT 135.580 -20.790 136.050 -19.870 ;
        RECT 142.330 -20.350 142.800 -19.420 ;
        RECT 149.080 -20.790 149.550 -19.870 ;
        RECT 155.830 -20.350 156.300 -19.420 ;
        RECT 162.580 -20.790 163.050 -19.870 ;
        RECT 169.330 -20.350 169.800 -19.420 ;
        RECT 176.080 -20.790 176.550 -19.870 ;
        RECT 182.830 -20.350 183.300 -19.420 ;
        RECT 189.580 -20.790 190.050 -19.870 ;
        RECT 196.330 -20.350 196.800 -19.420 ;
        RECT 203.080 -20.790 203.550 -19.870 ;
        RECT 209.830 -20.350 210.300 -19.420 ;
        RECT 216.580 -20.340 217.040 -19.870 ;
        RECT 216.580 -20.350 217.050 -20.340 ;
        RECT 216.590 -20.790 217.050 -20.350 ;
      LAYER via ;
        RECT 0.680 -20.200 0.950 -19.930 ;
        RECT 7.430 -20.250 7.700 -19.980 ;
        RECT 14.180 -20.200 14.450 -19.930 ;
        RECT 20.930 -20.220 21.200 -19.950 ;
        RECT 27.680 -20.200 27.950 -19.930 ;
        RECT 34.430 -20.220 34.700 -19.950 ;
        RECT 41.180 -20.200 41.450 -19.930 ;
        RECT 47.930 -20.250 48.200 -19.980 ;
        RECT 54.680 -20.200 54.950 -19.930 ;
        RECT 61.430 -20.250 61.700 -19.980 ;
        RECT 68.180 -20.200 68.450 -19.930 ;
        RECT 74.930 -20.220 75.200 -19.950 ;
        RECT 81.680 -20.200 81.950 -19.930 ;
        RECT 88.430 -20.220 88.700 -19.950 ;
        RECT 95.180 -20.200 95.450 -19.930 ;
        RECT 101.930 -20.250 102.200 -19.980 ;
        RECT 108.680 -20.200 108.950 -19.930 ;
        RECT 115.430 -20.250 115.700 -19.980 ;
        RECT 122.180 -20.200 122.450 -19.930 ;
        RECT 128.930 -20.220 129.200 -19.950 ;
        RECT 135.680 -20.200 135.950 -19.930 ;
        RECT 142.430 -20.220 142.700 -19.950 ;
        RECT 149.180 -20.200 149.450 -19.930 ;
        RECT 155.930 -20.250 156.200 -19.980 ;
        RECT 162.680 -20.200 162.950 -19.930 ;
        RECT 169.430 -20.250 169.700 -19.980 ;
        RECT 176.180 -20.200 176.450 -19.930 ;
        RECT 182.930 -20.220 183.200 -19.950 ;
        RECT 189.680 -20.200 189.950 -19.930 ;
        RECT 196.430 -20.220 196.700 -19.950 ;
        RECT 203.180 -20.200 203.450 -19.930 ;
        RECT 209.930 -20.250 210.200 -19.980 ;
        RECT 216.680 -20.200 216.950 -19.930 ;
      LAYER met2 ;
        RECT 0.580 -19.840 1.060 -19.830 ;
        RECT 14.040 -19.840 41.590 -19.830 ;
        RECT 68.040 -19.840 95.590 -19.830 ;
        RECT 108.570 -19.840 109.060 -19.830 ;
        RECT 122.040 -19.840 149.590 -19.830 ;
        RECT 176.040 -19.840 203.590 -19.830 ;
        RECT 216.570 -19.840 217.050 -19.830 ;
        RECT 0.580 -20.340 217.050 -19.840 ;
        RECT 0.590 -20.350 217.040 -20.340 ;
        RECT 0.590 -20.360 14.590 -20.350 ;
        RECT 41.040 -20.360 68.590 -20.350 ;
        RECT 95.040 -20.360 122.590 -20.350 ;
        RECT 149.040 -20.360 176.590 -20.350 ;
        RECT 203.040 -20.360 217.040 -20.350 ;
    END
  END WL20
  PIN WL21
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER li1 ;
        RECT 0.590 -21.680 1.040 -21.240 ;
        RECT 14.090 -21.680 14.540 -21.240 ;
        RECT 27.590 -21.680 28.040 -21.240 ;
        RECT 41.090 -21.680 41.540 -21.240 ;
        RECT 54.590 -21.680 55.040 -21.240 ;
        RECT 68.090 -21.680 68.540 -21.240 ;
        RECT 81.590 -21.680 82.040 -21.240 ;
        RECT 95.090 -21.680 95.540 -21.240 ;
        RECT 108.590 -21.680 109.040 -21.240 ;
        RECT 122.090 -21.680 122.540 -21.240 ;
        RECT 135.590 -21.680 136.040 -21.240 ;
        RECT 149.090 -21.680 149.540 -21.240 ;
        RECT 162.590 -21.680 163.040 -21.240 ;
        RECT 176.090 -21.680 176.540 -21.240 ;
        RECT 189.590 -21.680 190.040 -21.240 ;
        RECT 203.090 -21.680 203.540 -21.240 ;
        RECT 216.590 -21.680 217.040 -21.240 ;
        RECT 7.340 -22.600 7.790 -22.150 ;
        RECT 20.840 -22.600 21.290 -22.150 ;
        RECT 34.340 -22.600 34.790 -22.150 ;
        RECT 47.840 -22.600 48.290 -22.150 ;
        RECT 61.340 -22.600 61.790 -22.150 ;
        RECT 74.840 -22.600 75.290 -22.150 ;
        RECT 88.340 -22.600 88.790 -22.150 ;
        RECT 101.840 -22.600 102.290 -22.150 ;
        RECT 115.340 -22.600 115.790 -22.150 ;
        RECT 128.840 -22.600 129.290 -22.150 ;
        RECT 142.340 -22.600 142.790 -22.150 ;
        RECT 155.840 -22.600 156.290 -22.150 ;
        RECT 169.340 -22.600 169.790 -22.150 ;
        RECT 182.840 -22.600 183.290 -22.150 ;
        RECT 196.340 -22.600 196.790 -22.150 ;
        RECT 209.840 -22.600 210.290 -22.150 ;
      LAYER mcon ;
        RECT 0.680 -21.600 0.950 -21.330 ;
        RECT 14.180 -21.600 14.450 -21.330 ;
        RECT 27.680 -21.600 27.950 -21.330 ;
        RECT 41.180 -21.600 41.450 -21.330 ;
        RECT 54.680 -21.600 54.950 -21.330 ;
        RECT 68.180 -21.600 68.450 -21.330 ;
        RECT 81.680 -21.600 81.950 -21.330 ;
        RECT 95.180 -21.600 95.450 -21.330 ;
        RECT 108.680 -21.600 108.950 -21.330 ;
        RECT 122.180 -21.600 122.450 -21.330 ;
        RECT 135.680 -21.600 135.950 -21.330 ;
        RECT 149.180 -21.600 149.450 -21.330 ;
        RECT 162.680 -21.600 162.950 -21.330 ;
        RECT 176.180 -21.600 176.450 -21.330 ;
        RECT 189.680 -21.600 189.950 -21.330 ;
        RECT 203.180 -21.600 203.450 -21.330 ;
        RECT 216.680 -21.600 216.950 -21.330 ;
        RECT 7.440 -22.500 7.690 -22.250 ;
        RECT 20.940 -22.500 21.190 -22.250 ;
        RECT 34.440 -22.500 34.690 -22.250 ;
        RECT 47.940 -22.500 48.190 -22.250 ;
        RECT 61.440 -22.500 61.690 -22.250 ;
        RECT 74.940 -22.500 75.190 -22.250 ;
        RECT 88.440 -22.500 88.690 -22.250 ;
        RECT 101.940 -22.500 102.190 -22.250 ;
        RECT 115.440 -22.500 115.690 -22.250 ;
        RECT 128.940 -22.500 129.190 -22.250 ;
        RECT 142.440 -22.500 142.690 -22.250 ;
        RECT 155.940 -22.500 156.190 -22.250 ;
        RECT 169.440 -22.500 169.690 -22.250 ;
        RECT 182.940 -22.500 183.190 -22.250 ;
        RECT 196.440 -22.500 196.690 -22.250 ;
        RECT 209.940 -22.500 210.190 -22.250 ;
      LAYER met1 ;
        RECT 0.580 -21.680 1.040 -21.240 ;
        RECT 0.580 -21.690 1.050 -21.680 ;
        RECT 0.590 -22.160 1.050 -21.690 ;
        RECT 7.330 -22.610 7.800 -21.680 ;
        RECT 14.080 -22.160 14.550 -21.240 ;
        RECT 20.830 -22.610 21.300 -21.680 ;
        RECT 27.580 -22.160 28.050 -21.240 ;
        RECT 34.330 -22.610 34.800 -21.680 ;
        RECT 41.080 -22.160 41.550 -21.240 ;
        RECT 47.830 -22.610 48.300 -21.680 ;
        RECT 54.580 -22.160 55.050 -21.240 ;
        RECT 61.330 -22.610 61.800 -21.680 ;
        RECT 68.080 -22.160 68.550 -21.240 ;
        RECT 74.830 -22.610 75.300 -21.680 ;
        RECT 81.580 -22.160 82.050 -21.240 ;
        RECT 88.330 -22.610 88.800 -21.680 ;
        RECT 95.080 -22.160 95.550 -21.240 ;
        RECT 101.830 -22.610 102.300 -21.680 ;
        RECT 108.580 -22.160 109.050 -21.240 ;
        RECT 115.330 -22.610 115.800 -21.680 ;
        RECT 122.080 -22.160 122.550 -21.240 ;
        RECT 128.830 -22.610 129.300 -21.680 ;
        RECT 135.580 -22.160 136.050 -21.240 ;
        RECT 142.330 -22.610 142.800 -21.680 ;
        RECT 149.080 -22.160 149.550 -21.240 ;
        RECT 155.830 -22.610 156.300 -21.680 ;
        RECT 162.580 -22.160 163.050 -21.240 ;
        RECT 169.330 -22.610 169.800 -21.680 ;
        RECT 176.080 -22.160 176.550 -21.240 ;
        RECT 182.830 -22.610 183.300 -21.680 ;
        RECT 189.580 -22.160 190.050 -21.240 ;
        RECT 196.330 -22.610 196.800 -21.680 ;
        RECT 203.080 -22.160 203.550 -21.240 ;
        RECT 216.590 -21.680 217.050 -21.240 ;
        RECT 209.830 -22.610 210.300 -21.680 ;
        RECT 216.580 -21.690 217.050 -21.680 ;
        RECT 216.580 -22.160 217.040 -21.690 ;
      LAYER via ;
        RECT 0.680 -22.100 0.950 -21.830 ;
        RECT 7.430 -22.080 7.700 -21.810 ;
        RECT 14.180 -22.100 14.450 -21.830 ;
        RECT 20.930 -22.050 21.200 -21.780 ;
        RECT 27.680 -22.100 27.950 -21.830 ;
        RECT 34.430 -22.050 34.700 -21.780 ;
        RECT 41.180 -22.100 41.450 -21.830 ;
        RECT 47.930 -22.080 48.200 -21.810 ;
        RECT 54.680 -22.100 54.950 -21.830 ;
        RECT 61.430 -22.080 61.700 -21.810 ;
        RECT 68.180 -22.100 68.450 -21.830 ;
        RECT 74.930 -22.050 75.200 -21.780 ;
        RECT 81.680 -22.100 81.950 -21.830 ;
        RECT 88.430 -22.050 88.700 -21.780 ;
        RECT 95.180 -22.100 95.450 -21.830 ;
        RECT 101.930 -22.080 102.200 -21.810 ;
        RECT 108.680 -22.100 108.950 -21.830 ;
        RECT 115.430 -22.080 115.700 -21.810 ;
        RECT 122.180 -22.100 122.450 -21.830 ;
        RECT 128.930 -22.050 129.200 -21.780 ;
        RECT 135.680 -22.100 135.950 -21.830 ;
        RECT 142.430 -22.050 142.700 -21.780 ;
        RECT 149.180 -22.100 149.450 -21.830 ;
        RECT 155.930 -22.080 156.200 -21.810 ;
        RECT 162.680 -22.100 162.950 -21.830 ;
        RECT 169.430 -22.080 169.700 -21.810 ;
        RECT 176.180 -22.100 176.450 -21.830 ;
        RECT 182.930 -22.050 183.200 -21.780 ;
        RECT 189.680 -22.100 189.950 -21.830 ;
        RECT 196.430 -22.050 196.700 -21.780 ;
        RECT 203.180 -22.100 203.450 -21.830 ;
        RECT 209.930 -22.080 210.200 -21.810 ;
        RECT 216.680 -22.100 216.950 -21.830 ;
      LAYER met2 ;
        RECT 14.040 -21.680 41.590 -21.670 ;
        RECT 68.040 -21.680 95.590 -21.670 ;
        RECT 122.040 -21.680 149.590 -21.670 ;
        RECT 176.040 -21.680 203.590 -21.670 ;
        RECT 0.590 -21.690 217.040 -21.680 ;
        RECT 0.580 -22.190 217.050 -21.690 ;
        RECT 0.580 -22.200 14.590 -22.190 ;
        RECT 41.040 -22.200 68.590 -22.190 ;
        RECT 95.040 -22.200 122.590 -22.190 ;
        RECT 149.040 -22.200 176.590 -22.190 ;
        RECT 203.040 -22.200 217.050 -22.190 ;
        RECT 0.580 -22.210 1.060 -22.200 ;
        RECT 108.570 -22.210 109.060 -22.200 ;
        RECT 216.570 -22.210 217.050 -22.200 ;
    END
  END WL21
  PIN WL22
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER li1 ;
        RECT 7.340 -23.490 7.790 -23.040 ;
        RECT 20.840 -23.490 21.290 -23.040 ;
        RECT 34.340 -23.490 34.790 -23.040 ;
        RECT 47.840 -23.490 48.290 -23.040 ;
        RECT 61.340 -23.490 61.790 -23.040 ;
        RECT 74.840 -23.490 75.290 -23.040 ;
        RECT 88.340 -23.490 88.790 -23.040 ;
        RECT 101.840 -23.490 102.290 -23.040 ;
        RECT 115.340 -23.490 115.790 -23.040 ;
        RECT 128.840 -23.490 129.290 -23.040 ;
        RECT 142.340 -23.490 142.790 -23.040 ;
        RECT 155.840 -23.490 156.290 -23.040 ;
        RECT 169.340 -23.490 169.790 -23.040 ;
        RECT 182.840 -23.490 183.290 -23.040 ;
        RECT 196.340 -23.490 196.790 -23.040 ;
        RECT 209.840 -23.490 210.290 -23.040 ;
        RECT 0.590 -24.400 1.040 -23.960 ;
        RECT 14.090 -24.400 14.540 -23.960 ;
        RECT 27.590 -24.400 28.040 -23.960 ;
        RECT 41.090 -24.400 41.540 -23.960 ;
        RECT 54.590 -24.400 55.040 -23.960 ;
        RECT 68.090 -24.400 68.540 -23.960 ;
        RECT 81.590 -24.400 82.040 -23.960 ;
        RECT 95.090 -24.400 95.540 -23.960 ;
        RECT 108.590 -24.400 109.040 -23.960 ;
        RECT 122.090 -24.400 122.540 -23.960 ;
        RECT 135.590 -24.400 136.040 -23.960 ;
        RECT 149.090 -24.400 149.540 -23.960 ;
        RECT 162.590 -24.400 163.040 -23.960 ;
        RECT 176.090 -24.400 176.540 -23.960 ;
        RECT 189.590 -24.400 190.040 -23.960 ;
        RECT 203.090 -24.400 203.540 -23.960 ;
        RECT 216.590 -24.400 217.040 -23.960 ;
      LAYER mcon ;
        RECT 7.440 -23.390 7.690 -23.140 ;
        RECT 20.940 -23.390 21.190 -23.140 ;
        RECT 34.440 -23.390 34.690 -23.140 ;
        RECT 47.940 -23.390 48.190 -23.140 ;
        RECT 61.440 -23.390 61.690 -23.140 ;
        RECT 74.940 -23.390 75.190 -23.140 ;
        RECT 88.440 -23.390 88.690 -23.140 ;
        RECT 101.940 -23.390 102.190 -23.140 ;
        RECT 115.440 -23.390 115.690 -23.140 ;
        RECT 128.940 -23.390 129.190 -23.140 ;
        RECT 142.440 -23.390 142.690 -23.140 ;
        RECT 155.940 -23.390 156.190 -23.140 ;
        RECT 169.440 -23.390 169.690 -23.140 ;
        RECT 182.940 -23.390 183.190 -23.140 ;
        RECT 196.440 -23.390 196.690 -23.140 ;
        RECT 209.940 -23.390 210.190 -23.140 ;
        RECT 0.680 -24.310 0.950 -24.040 ;
        RECT 14.180 -24.310 14.450 -24.040 ;
        RECT 27.680 -24.310 27.950 -24.040 ;
        RECT 41.180 -24.310 41.450 -24.040 ;
        RECT 54.680 -24.310 54.950 -24.040 ;
        RECT 68.180 -24.310 68.450 -24.040 ;
        RECT 81.680 -24.310 81.950 -24.040 ;
        RECT 95.180 -24.310 95.450 -24.040 ;
        RECT 108.680 -24.310 108.950 -24.040 ;
        RECT 122.180 -24.310 122.450 -24.040 ;
        RECT 135.680 -24.310 135.950 -24.040 ;
        RECT 149.180 -24.310 149.450 -24.040 ;
        RECT 162.680 -24.310 162.950 -24.040 ;
        RECT 176.180 -24.310 176.450 -24.040 ;
        RECT 189.680 -24.310 189.950 -24.040 ;
        RECT 203.180 -24.310 203.450 -24.040 ;
        RECT 216.680 -24.310 216.950 -24.040 ;
      LAYER met1 ;
        RECT 0.590 -23.950 1.050 -23.480 ;
        RECT 0.580 -23.960 1.050 -23.950 ;
        RECT 7.330 -23.960 7.800 -23.030 ;
        RECT 0.580 -24.400 1.040 -23.960 ;
        RECT 14.080 -24.400 14.550 -23.480 ;
        RECT 20.830 -23.960 21.300 -23.030 ;
        RECT 27.580 -24.400 28.050 -23.480 ;
        RECT 34.330 -23.960 34.800 -23.030 ;
        RECT 41.080 -24.400 41.550 -23.480 ;
        RECT 47.830 -23.960 48.300 -23.030 ;
        RECT 54.580 -24.400 55.050 -23.480 ;
        RECT 61.330 -23.960 61.800 -23.030 ;
        RECT 68.080 -24.400 68.550 -23.480 ;
        RECT 74.830 -23.960 75.300 -23.030 ;
        RECT 81.580 -24.400 82.050 -23.480 ;
        RECT 88.330 -23.960 88.800 -23.030 ;
        RECT 95.080 -24.400 95.550 -23.480 ;
        RECT 101.830 -23.960 102.300 -23.030 ;
        RECT 108.580 -24.400 109.050 -23.480 ;
        RECT 115.330 -23.960 115.800 -23.030 ;
        RECT 122.080 -24.400 122.550 -23.480 ;
        RECT 128.830 -23.960 129.300 -23.030 ;
        RECT 135.580 -24.400 136.050 -23.480 ;
        RECT 142.330 -23.960 142.800 -23.030 ;
        RECT 149.080 -24.400 149.550 -23.480 ;
        RECT 155.830 -23.960 156.300 -23.030 ;
        RECT 162.580 -24.400 163.050 -23.480 ;
        RECT 169.330 -23.960 169.800 -23.030 ;
        RECT 176.080 -24.400 176.550 -23.480 ;
        RECT 182.830 -23.960 183.300 -23.030 ;
        RECT 189.580 -24.400 190.050 -23.480 ;
        RECT 196.330 -23.960 196.800 -23.030 ;
        RECT 203.080 -24.400 203.550 -23.480 ;
        RECT 209.830 -23.960 210.300 -23.030 ;
        RECT 216.580 -23.950 217.040 -23.480 ;
        RECT 216.580 -23.960 217.050 -23.950 ;
        RECT 216.590 -24.400 217.050 -23.960 ;
      LAYER via ;
        RECT 0.680 -23.810 0.950 -23.540 ;
        RECT 7.430 -23.860 7.700 -23.590 ;
        RECT 14.180 -23.810 14.450 -23.540 ;
        RECT 20.930 -23.860 21.200 -23.590 ;
        RECT 27.680 -23.810 27.950 -23.540 ;
        RECT 34.430 -23.860 34.700 -23.590 ;
        RECT 41.180 -23.810 41.450 -23.540 ;
        RECT 47.930 -23.860 48.200 -23.590 ;
        RECT 54.680 -23.810 54.950 -23.540 ;
        RECT 61.430 -23.860 61.700 -23.590 ;
        RECT 68.180 -23.810 68.450 -23.540 ;
        RECT 74.930 -23.860 75.200 -23.590 ;
        RECT 81.680 -23.810 81.950 -23.540 ;
        RECT 88.430 -23.860 88.700 -23.590 ;
        RECT 95.180 -23.810 95.450 -23.540 ;
        RECT 101.930 -23.860 102.200 -23.590 ;
        RECT 108.680 -23.810 108.950 -23.540 ;
        RECT 115.430 -23.860 115.700 -23.590 ;
        RECT 122.180 -23.810 122.450 -23.540 ;
        RECT 128.930 -23.860 129.200 -23.590 ;
        RECT 135.680 -23.810 135.950 -23.540 ;
        RECT 142.430 -23.860 142.700 -23.590 ;
        RECT 149.180 -23.810 149.450 -23.540 ;
        RECT 155.930 -23.860 156.200 -23.590 ;
        RECT 162.680 -23.810 162.950 -23.540 ;
        RECT 169.430 -23.860 169.700 -23.590 ;
        RECT 176.180 -23.810 176.450 -23.540 ;
        RECT 182.930 -23.860 183.200 -23.590 ;
        RECT 189.680 -23.810 189.950 -23.540 ;
        RECT 196.430 -23.860 196.700 -23.590 ;
        RECT 203.180 -23.810 203.450 -23.540 ;
        RECT 209.930 -23.860 210.200 -23.590 ;
        RECT 216.680 -23.810 216.950 -23.540 ;
      LAYER met2 ;
        RECT 0.590 -23.970 217.040 -23.450 ;
    END
  END WL22
  PIN WL23
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER li1 ;
        RECT 0.590 -25.290 1.040 -24.850 ;
        RECT 14.090 -25.290 14.540 -24.850 ;
        RECT 27.590 -25.290 28.040 -24.850 ;
        RECT 41.090 -25.290 41.540 -24.850 ;
        RECT 54.590 -25.290 55.040 -24.850 ;
        RECT 68.090 -25.290 68.540 -24.850 ;
        RECT 81.590 -25.290 82.040 -24.850 ;
        RECT 95.090 -25.290 95.540 -24.850 ;
        RECT 108.590 -25.290 109.040 -24.850 ;
        RECT 122.090 -25.290 122.540 -24.850 ;
        RECT 135.590 -25.290 136.040 -24.850 ;
        RECT 149.090 -25.290 149.540 -24.850 ;
        RECT 162.590 -25.290 163.040 -24.850 ;
        RECT 176.090 -25.290 176.540 -24.850 ;
        RECT 189.590 -25.290 190.040 -24.850 ;
        RECT 203.090 -25.290 203.540 -24.850 ;
        RECT 216.590 -25.290 217.040 -24.850 ;
        RECT 7.340 -26.210 7.790 -25.760 ;
        RECT 20.840 -26.210 21.290 -25.760 ;
        RECT 34.340 -26.210 34.790 -25.760 ;
        RECT 47.840 -26.210 48.290 -25.760 ;
        RECT 61.340 -26.210 61.790 -25.760 ;
        RECT 74.840 -26.210 75.290 -25.760 ;
        RECT 88.340 -26.210 88.790 -25.760 ;
        RECT 101.840 -26.210 102.290 -25.760 ;
        RECT 115.340 -26.210 115.790 -25.760 ;
        RECT 128.840 -26.210 129.290 -25.760 ;
        RECT 142.340 -26.210 142.790 -25.760 ;
        RECT 155.840 -26.210 156.290 -25.760 ;
        RECT 169.340 -26.210 169.790 -25.760 ;
        RECT 182.840 -26.210 183.290 -25.760 ;
        RECT 196.340 -26.210 196.790 -25.760 ;
        RECT 209.840 -26.210 210.290 -25.760 ;
      LAYER mcon ;
        RECT 0.680 -25.210 0.950 -24.940 ;
        RECT 14.180 -25.210 14.450 -24.940 ;
        RECT 27.680 -25.210 27.950 -24.940 ;
        RECT 41.180 -25.210 41.450 -24.940 ;
        RECT 54.680 -25.210 54.950 -24.940 ;
        RECT 68.180 -25.210 68.450 -24.940 ;
        RECT 81.680 -25.210 81.950 -24.940 ;
        RECT 95.180 -25.210 95.450 -24.940 ;
        RECT 108.680 -25.210 108.950 -24.940 ;
        RECT 122.180 -25.210 122.450 -24.940 ;
        RECT 135.680 -25.210 135.950 -24.940 ;
        RECT 149.180 -25.210 149.450 -24.940 ;
        RECT 162.680 -25.210 162.950 -24.940 ;
        RECT 176.180 -25.210 176.450 -24.940 ;
        RECT 189.680 -25.210 189.950 -24.940 ;
        RECT 203.180 -25.210 203.450 -24.940 ;
        RECT 216.680 -25.210 216.950 -24.940 ;
        RECT 7.440 -26.110 7.690 -25.860 ;
        RECT 20.940 -26.110 21.190 -25.860 ;
        RECT 34.440 -26.110 34.690 -25.860 ;
        RECT 47.940 -26.110 48.190 -25.860 ;
        RECT 61.440 -26.110 61.690 -25.860 ;
        RECT 74.940 -26.110 75.190 -25.860 ;
        RECT 88.440 -26.110 88.690 -25.860 ;
        RECT 101.940 -26.110 102.190 -25.860 ;
        RECT 115.440 -26.110 115.690 -25.860 ;
        RECT 128.940 -26.110 129.190 -25.860 ;
        RECT 142.440 -26.110 142.690 -25.860 ;
        RECT 155.940 -26.110 156.190 -25.860 ;
        RECT 169.440 -26.110 169.690 -25.860 ;
        RECT 182.940 -26.110 183.190 -25.860 ;
        RECT 196.440 -26.110 196.690 -25.860 ;
        RECT 209.940 -26.110 210.190 -25.860 ;
      LAYER met1 ;
        RECT 0.580 -25.290 1.040 -24.850 ;
        RECT 0.580 -25.300 1.050 -25.290 ;
        RECT 0.590 -25.770 1.050 -25.300 ;
        RECT 7.330 -26.220 7.800 -25.290 ;
        RECT 14.080 -25.770 14.550 -24.850 ;
        RECT 20.830 -26.220 21.300 -25.290 ;
        RECT 27.580 -25.770 28.050 -24.850 ;
        RECT 34.330 -26.220 34.800 -25.290 ;
        RECT 41.080 -25.770 41.550 -24.850 ;
        RECT 47.830 -26.220 48.300 -25.290 ;
        RECT 54.580 -25.770 55.050 -24.850 ;
        RECT 61.330 -26.220 61.800 -25.290 ;
        RECT 68.080 -25.770 68.550 -24.850 ;
        RECT 74.830 -26.220 75.300 -25.290 ;
        RECT 81.580 -25.770 82.050 -24.850 ;
        RECT 88.330 -26.220 88.800 -25.290 ;
        RECT 95.080 -25.770 95.550 -24.850 ;
        RECT 101.830 -26.220 102.300 -25.290 ;
        RECT 108.580 -25.770 109.050 -24.850 ;
        RECT 115.330 -26.220 115.800 -25.290 ;
        RECT 122.080 -25.770 122.550 -24.850 ;
        RECT 128.830 -26.220 129.300 -25.290 ;
        RECT 135.580 -25.770 136.050 -24.850 ;
        RECT 142.330 -26.220 142.800 -25.290 ;
        RECT 149.080 -25.770 149.550 -24.850 ;
        RECT 155.830 -26.220 156.300 -25.290 ;
        RECT 162.580 -25.770 163.050 -24.850 ;
        RECT 169.330 -26.220 169.800 -25.290 ;
        RECT 176.080 -25.770 176.550 -24.850 ;
        RECT 182.830 -26.220 183.300 -25.290 ;
        RECT 189.580 -25.770 190.050 -24.850 ;
        RECT 196.330 -26.220 196.800 -25.290 ;
        RECT 203.080 -25.770 203.550 -24.850 ;
        RECT 216.590 -25.290 217.050 -24.850 ;
        RECT 209.830 -26.220 210.300 -25.290 ;
        RECT 216.580 -25.300 217.050 -25.290 ;
        RECT 216.580 -25.770 217.040 -25.300 ;
      LAYER via ;
        RECT 0.680 -25.710 0.950 -25.440 ;
        RECT 7.430 -25.690 7.700 -25.420 ;
        RECT 14.180 -25.710 14.450 -25.440 ;
        RECT 20.930 -25.690 21.200 -25.420 ;
        RECT 27.680 -25.710 27.950 -25.440 ;
        RECT 34.430 -25.690 34.700 -25.420 ;
        RECT 41.180 -25.710 41.450 -25.440 ;
        RECT 47.930 -25.690 48.200 -25.420 ;
        RECT 54.680 -25.710 54.950 -25.440 ;
        RECT 61.430 -25.690 61.700 -25.420 ;
        RECT 68.180 -25.710 68.450 -25.440 ;
        RECT 74.930 -25.690 75.200 -25.420 ;
        RECT 81.680 -25.710 81.950 -25.440 ;
        RECT 88.430 -25.690 88.700 -25.420 ;
        RECT 95.180 -25.710 95.450 -25.440 ;
        RECT 101.930 -25.690 102.200 -25.420 ;
        RECT 108.680 -25.710 108.950 -25.440 ;
        RECT 115.430 -25.690 115.700 -25.420 ;
        RECT 122.180 -25.710 122.450 -25.440 ;
        RECT 128.930 -25.690 129.200 -25.420 ;
        RECT 135.680 -25.710 135.950 -25.440 ;
        RECT 142.430 -25.690 142.700 -25.420 ;
        RECT 149.180 -25.710 149.450 -25.440 ;
        RECT 155.930 -25.690 156.200 -25.420 ;
        RECT 162.680 -25.710 162.950 -25.440 ;
        RECT 169.430 -25.690 169.700 -25.420 ;
        RECT 176.180 -25.710 176.450 -25.440 ;
        RECT 182.930 -25.690 183.200 -25.420 ;
        RECT 189.680 -25.710 189.950 -25.440 ;
        RECT 196.430 -25.690 196.700 -25.420 ;
        RECT 203.180 -25.710 203.450 -25.440 ;
        RECT 209.930 -25.690 210.200 -25.420 ;
        RECT 216.680 -25.710 216.950 -25.440 ;
      LAYER met2 ;
        RECT 0.590 -25.310 217.040 -25.290 ;
        RECT 0.580 -25.810 217.050 -25.310 ;
        RECT 0.580 -25.820 1.060 -25.810 ;
        RECT 108.570 -25.820 109.060 -25.810 ;
        RECT 216.570 -25.820 217.050 -25.810 ;
    END
  END WL23
  PIN WL24
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER li1 ;
        RECT 7.340 -27.100 7.790 -26.650 ;
        RECT 20.840 -27.100 21.290 -26.650 ;
        RECT 34.340 -27.100 34.790 -26.650 ;
        RECT 47.840 -27.100 48.290 -26.650 ;
        RECT 61.340 -27.100 61.790 -26.650 ;
        RECT 74.840 -27.100 75.290 -26.650 ;
        RECT 88.340 -27.100 88.790 -26.650 ;
        RECT 101.840 -27.100 102.290 -26.650 ;
        RECT 115.340 -27.100 115.790 -26.650 ;
        RECT 128.840 -27.100 129.290 -26.650 ;
        RECT 142.340 -27.100 142.790 -26.650 ;
        RECT 155.840 -27.100 156.290 -26.650 ;
        RECT 169.340 -27.100 169.790 -26.650 ;
        RECT 182.840 -27.100 183.290 -26.650 ;
        RECT 196.340 -27.100 196.790 -26.650 ;
        RECT 209.840 -27.100 210.290 -26.650 ;
        RECT 0.590 -28.010 1.040 -27.570 ;
        RECT 14.090 -28.010 14.540 -27.570 ;
        RECT 27.590 -28.010 28.040 -27.570 ;
        RECT 41.090 -28.010 41.540 -27.570 ;
        RECT 54.590 -28.010 55.040 -27.570 ;
        RECT 68.090 -28.010 68.540 -27.570 ;
        RECT 81.590 -28.010 82.040 -27.570 ;
        RECT 95.090 -28.010 95.540 -27.570 ;
        RECT 108.590 -28.010 109.040 -27.570 ;
        RECT 122.090 -28.010 122.540 -27.570 ;
        RECT 135.590 -28.010 136.040 -27.570 ;
        RECT 149.090 -28.010 149.540 -27.570 ;
        RECT 162.590 -28.010 163.040 -27.570 ;
        RECT 176.090 -28.010 176.540 -27.570 ;
        RECT 189.590 -28.010 190.040 -27.570 ;
        RECT 203.090 -28.010 203.540 -27.570 ;
        RECT 216.590 -28.010 217.040 -27.570 ;
      LAYER mcon ;
        RECT 7.440 -27.000 7.690 -26.750 ;
        RECT 20.940 -27.000 21.190 -26.750 ;
        RECT 34.440 -27.000 34.690 -26.750 ;
        RECT 47.940 -27.000 48.190 -26.750 ;
        RECT 61.440 -27.000 61.690 -26.750 ;
        RECT 74.940 -27.000 75.190 -26.750 ;
        RECT 88.440 -27.000 88.690 -26.750 ;
        RECT 101.940 -27.000 102.190 -26.750 ;
        RECT 115.440 -27.000 115.690 -26.750 ;
        RECT 128.940 -27.000 129.190 -26.750 ;
        RECT 142.440 -27.000 142.690 -26.750 ;
        RECT 155.940 -27.000 156.190 -26.750 ;
        RECT 169.440 -27.000 169.690 -26.750 ;
        RECT 182.940 -27.000 183.190 -26.750 ;
        RECT 196.440 -27.000 196.690 -26.750 ;
        RECT 209.940 -27.000 210.190 -26.750 ;
        RECT 0.680 -27.920 0.950 -27.650 ;
        RECT 14.180 -27.920 14.450 -27.650 ;
        RECT 27.680 -27.920 27.950 -27.650 ;
        RECT 41.180 -27.920 41.450 -27.650 ;
        RECT 54.680 -27.920 54.950 -27.650 ;
        RECT 68.180 -27.920 68.450 -27.650 ;
        RECT 81.680 -27.920 81.950 -27.650 ;
        RECT 95.180 -27.920 95.450 -27.650 ;
        RECT 108.680 -27.920 108.950 -27.650 ;
        RECT 122.180 -27.920 122.450 -27.650 ;
        RECT 135.680 -27.920 135.950 -27.650 ;
        RECT 149.180 -27.920 149.450 -27.650 ;
        RECT 162.680 -27.920 162.950 -27.650 ;
        RECT 176.180 -27.920 176.450 -27.650 ;
        RECT 189.680 -27.920 189.950 -27.650 ;
        RECT 203.180 -27.920 203.450 -27.650 ;
        RECT 216.680 -27.920 216.950 -27.650 ;
      LAYER met1 ;
        RECT 0.590 -27.560 1.050 -27.090 ;
        RECT 0.580 -27.570 1.050 -27.560 ;
        RECT 7.330 -27.570 7.800 -26.640 ;
        RECT 0.580 -28.010 1.040 -27.570 ;
        RECT 14.080 -28.010 14.550 -27.090 ;
        RECT 20.830 -27.570 21.300 -26.640 ;
        RECT 27.580 -28.010 28.050 -27.090 ;
        RECT 34.330 -27.570 34.800 -26.640 ;
        RECT 41.080 -28.010 41.550 -27.090 ;
        RECT 47.830 -27.570 48.300 -26.640 ;
        RECT 54.580 -28.010 55.050 -27.090 ;
        RECT 61.330 -27.570 61.800 -26.640 ;
        RECT 68.080 -28.010 68.550 -27.090 ;
        RECT 74.830 -27.570 75.300 -26.640 ;
        RECT 81.580 -28.010 82.050 -27.090 ;
        RECT 88.330 -27.570 88.800 -26.640 ;
        RECT 95.080 -28.010 95.550 -27.090 ;
        RECT 101.830 -27.570 102.300 -26.640 ;
        RECT 108.580 -28.010 109.050 -27.090 ;
        RECT 115.330 -27.570 115.800 -26.640 ;
        RECT 122.080 -28.010 122.550 -27.090 ;
        RECT 128.830 -27.570 129.300 -26.640 ;
        RECT 135.580 -28.010 136.050 -27.090 ;
        RECT 142.330 -27.570 142.800 -26.640 ;
        RECT 149.080 -28.010 149.550 -27.090 ;
        RECT 155.830 -27.570 156.300 -26.640 ;
        RECT 162.580 -28.010 163.050 -27.090 ;
        RECT 169.330 -27.570 169.800 -26.640 ;
        RECT 176.080 -28.010 176.550 -27.090 ;
        RECT 182.830 -27.570 183.300 -26.640 ;
        RECT 189.580 -28.010 190.050 -27.090 ;
        RECT 196.330 -27.570 196.800 -26.640 ;
        RECT 203.080 -28.010 203.550 -27.090 ;
        RECT 209.830 -27.570 210.300 -26.640 ;
        RECT 216.580 -27.560 217.040 -27.090 ;
        RECT 216.580 -27.570 217.050 -27.560 ;
        RECT 216.590 -28.010 217.050 -27.570 ;
      LAYER via ;
        RECT 0.680 -27.420 0.950 -27.150 ;
        RECT 7.430 -27.440 7.700 -27.170 ;
        RECT 14.180 -27.420 14.450 -27.150 ;
        RECT 20.930 -27.440 21.200 -27.170 ;
        RECT 27.680 -27.420 27.950 -27.150 ;
        RECT 34.430 -27.440 34.700 -27.170 ;
        RECT 41.180 -27.420 41.450 -27.150 ;
        RECT 47.930 -27.440 48.200 -27.170 ;
        RECT 54.680 -27.420 54.950 -27.150 ;
        RECT 61.430 -27.440 61.700 -27.170 ;
        RECT 68.180 -27.420 68.450 -27.150 ;
        RECT 74.930 -27.440 75.200 -27.170 ;
        RECT 81.680 -27.420 81.950 -27.150 ;
        RECT 88.430 -27.440 88.700 -27.170 ;
        RECT 95.180 -27.420 95.450 -27.150 ;
        RECT 101.930 -27.440 102.200 -27.170 ;
        RECT 108.680 -27.420 108.950 -27.150 ;
        RECT 115.430 -27.440 115.700 -27.170 ;
        RECT 122.180 -27.420 122.450 -27.150 ;
        RECT 128.930 -27.440 129.200 -27.170 ;
        RECT 135.680 -27.420 135.950 -27.150 ;
        RECT 142.430 -27.440 142.700 -27.170 ;
        RECT 149.180 -27.420 149.450 -27.150 ;
        RECT 155.930 -27.440 156.200 -27.170 ;
        RECT 162.680 -27.420 162.950 -27.150 ;
        RECT 169.430 -27.440 169.700 -27.170 ;
        RECT 176.180 -27.420 176.450 -27.150 ;
        RECT 182.930 -27.440 183.200 -27.170 ;
        RECT 189.680 -27.420 189.950 -27.150 ;
        RECT 196.430 -27.440 196.700 -27.170 ;
        RECT 203.180 -27.420 203.450 -27.150 ;
        RECT 209.930 -27.440 210.200 -27.170 ;
        RECT 216.680 -27.420 216.950 -27.150 ;
      LAYER met2 ;
        RECT 0.580 -27.050 1.060 -27.040 ;
        RECT 108.570 -27.050 109.060 -27.040 ;
        RECT 216.570 -27.050 217.050 -27.040 ;
        RECT 0.580 -27.550 217.050 -27.050 ;
        RECT 0.590 -27.570 217.040 -27.550 ;
    END
  END WL24
  PIN WL25
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER li1 ;
        RECT 0.590 -28.900 1.040 -28.460 ;
        RECT 14.090 -28.900 14.540 -28.460 ;
        RECT 27.590 -28.900 28.040 -28.460 ;
        RECT 41.090 -28.900 41.540 -28.460 ;
        RECT 54.590 -28.900 55.040 -28.460 ;
        RECT 68.090 -28.900 68.540 -28.460 ;
        RECT 81.590 -28.900 82.040 -28.460 ;
        RECT 95.090 -28.900 95.540 -28.460 ;
        RECT 108.590 -28.900 109.040 -28.460 ;
        RECT 122.090 -28.900 122.540 -28.460 ;
        RECT 135.590 -28.900 136.040 -28.460 ;
        RECT 149.090 -28.900 149.540 -28.460 ;
        RECT 162.590 -28.900 163.040 -28.460 ;
        RECT 176.090 -28.900 176.540 -28.460 ;
        RECT 189.590 -28.900 190.040 -28.460 ;
        RECT 203.090 -28.900 203.540 -28.460 ;
        RECT 216.590 -28.900 217.040 -28.460 ;
        RECT 7.340 -29.820 7.790 -29.370 ;
        RECT 20.840 -29.820 21.290 -29.370 ;
        RECT 34.340 -29.820 34.790 -29.370 ;
        RECT 47.840 -29.820 48.290 -29.370 ;
        RECT 61.340 -29.820 61.790 -29.370 ;
        RECT 74.840 -29.820 75.290 -29.370 ;
        RECT 88.340 -29.820 88.790 -29.370 ;
        RECT 101.840 -29.820 102.290 -29.370 ;
        RECT 115.340 -29.820 115.790 -29.370 ;
        RECT 128.840 -29.820 129.290 -29.370 ;
        RECT 142.340 -29.820 142.790 -29.370 ;
        RECT 155.840 -29.820 156.290 -29.370 ;
        RECT 169.340 -29.820 169.790 -29.370 ;
        RECT 182.840 -29.820 183.290 -29.370 ;
        RECT 196.340 -29.820 196.790 -29.370 ;
        RECT 209.840 -29.820 210.290 -29.370 ;
      LAYER mcon ;
        RECT 0.680 -28.820 0.950 -28.550 ;
        RECT 14.180 -28.820 14.450 -28.550 ;
        RECT 27.680 -28.820 27.950 -28.550 ;
        RECT 41.180 -28.820 41.450 -28.550 ;
        RECT 54.680 -28.820 54.950 -28.550 ;
        RECT 68.180 -28.820 68.450 -28.550 ;
        RECT 81.680 -28.820 81.950 -28.550 ;
        RECT 95.180 -28.820 95.450 -28.550 ;
        RECT 108.680 -28.820 108.950 -28.550 ;
        RECT 122.180 -28.820 122.450 -28.550 ;
        RECT 135.680 -28.820 135.950 -28.550 ;
        RECT 149.180 -28.820 149.450 -28.550 ;
        RECT 162.680 -28.820 162.950 -28.550 ;
        RECT 176.180 -28.820 176.450 -28.550 ;
        RECT 189.680 -28.820 189.950 -28.550 ;
        RECT 203.180 -28.820 203.450 -28.550 ;
        RECT 216.680 -28.820 216.950 -28.550 ;
        RECT 7.440 -29.720 7.690 -29.470 ;
        RECT 20.940 -29.720 21.190 -29.470 ;
        RECT 34.440 -29.720 34.690 -29.470 ;
        RECT 47.940 -29.720 48.190 -29.470 ;
        RECT 61.440 -29.720 61.690 -29.470 ;
        RECT 74.940 -29.720 75.190 -29.470 ;
        RECT 88.440 -29.720 88.690 -29.470 ;
        RECT 101.940 -29.720 102.190 -29.470 ;
        RECT 115.440 -29.720 115.690 -29.470 ;
        RECT 128.940 -29.720 129.190 -29.470 ;
        RECT 142.440 -29.720 142.690 -29.470 ;
        RECT 155.940 -29.720 156.190 -29.470 ;
        RECT 169.440 -29.720 169.690 -29.470 ;
        RECT 182.940 -29.720 183.190 -29.470 ;
        RECT 196.440 -29.720 196.690 -29.470 ;
        RECT 209.940 -29.720 210.190 -29.470 ;
      LAYER met1 ;
        RECT 0.580 -28.900 1.040 -28.460 ;
        RECT 0.580 -28.910 1.050 -28.900 ;
        RECT 0.590 -29.380 1.050 -28.910 ;
        RECT 7.330 -29.830 7.800 -28.900 ;
        RECT 14.080 -29.380 14.550 -28.460 ;
        RECT 20.830 -29.830 21.300 -28.900 ;
        RECT 27.580 -29.380 28.050 -28.460 ;
        RECT 34.330 -29.830 34.800 -28.900 ;
        RECT 41.080 -29.380 41.550 -28.460 ;
        RECT 47.830 -29.830 48.300 -28.900 ;
        RECT 54.580 -29.380 55.050 -28.460 ;
        RECT 61.330 -29.830 61.800 -28.900 ;
        RECT 68.080 -29.380 68.550 -28.460 ;
        RECT 74.830 -29.830 75.300 -28.900 ;
        RECT 81.580 -29.380 82.050 -28.460 ;
        RECT 88.330 -29.830 88.800 -28.900 ;
        RECT 95.080 -29.380 95.550 -28.460 ;
        RECT 101.830 -29.830 102.300 -28.900 ;
        RECT 108.580 -29.380 109.050 -28.460 ;
        RECT 115.330 -29.830 115.800 -28.900 ;
        RECT 122.080 -29.380 122.550 -28.460 ;
        RECT 128.830 -29.830 129.300 -28.900 ;
        RECT 135.580 -29.380 136.050 -28.460 ;
        RECT 142.330 -29.830 142.800 -28.900 ;
        RECT 149.080 -29.380 149.550 -28.460 ;
        RECT 155.830 -29.830 156.300 -28.900 ;
        RECT 162.580 -29.380 163.050 -28.460 ;
        RECT 169.330 -29.830 169.800 -28.900 ;
        RECT 176.080 -29.380 176.550 -28.460 ;
        RECT 182.830 -29.830 183.300 -28.900 ;
        RECT 189.580 -29.380 190.050 -28.460 ;
        RECT 196.330 -29.830 196.800 -28.900 ;
        RECT 203.080 -29.380 203.550 -28.460 ;
        RECT 216.590 -28.900 217.050 -28.460 ;
        RECT 209.830 -29.830 210.300 -28.900 ;
        RECT 216.580 -28.910 217.050 -28.900 ;
        RECT 216.580 -29.380 217.040 -28.910 ;
      LAYER via ;
        RECT 0.680 -29.320 0.950 -29.050 ;
        RECT 7.430 -29.270 7.700 -29.000 ;
        RECT 14.180 -29.320 14.450 -29.050 ;
        RECT 20.930 -29.270 21.200 -29.000 ;
        RECT 27.680 -29.320 27.950 -29.050 ;
        RECT 34.430 -29.270 34.700 -29.000 ;
        RECT 41.180 -29.320 41.450 -29.050 ;
        RECT 47.930 -29.270 48.200 -29.000 ;
        RECT 54.680 -29.320 54.950 -29.050 ;
        RECT 61.430 -29.270 61.700 -29.000 ;
        RECT 68.180 -29.320 68.450 -29.050 ;
        RECT 74.930 -29.270 75.200 -29.000 ;
        RECT 81.680 -29.320 81.950 -29.050 ;
        RECT 88.430 -29.270 88.700 -29.000 ;
        RECT 95.180 -29.320 95.450 -29.050 ;
        RECT 101.930 -29.270 102.200 -29.000 ;
        RECT 108.680 -29.320 108.950 -29.050 ;
        RECT 115.430 -29.270 115.700 -29.000 ;
        RECT 122.180 -29.320 122.450 -29.050 ;
        RECT 128.930 -29.270 129.200 -29.000 ;
        RECT 135.680 -29.320 135.950 -29.050 ;
        RECT 142.430 -29.270 142.700 -29.000 ;
        RECT 149.180 -29.320 149.450 -29.050 ;
        RECT 155.930 -29.270 156.200 -29.000 ;
        RECT 162.680 -29.320 162.950 -29.050 ;
        RECT 169.430 -29.270 169.700 -29.000 ;
        RECT 176.180 -29.320 176.450 -29.050 ;
        RECT 182.930 -29.270 183.200 -29.000 ;
        RECT 189.680 -29.320 189.950 -29.050 ;
        RECT 196.430 -29.270 196.700 -29.000 ;
        RECT 203.180 -29.320 203.450 -29.050 ;
        RECT 209.930 -29.270 210.200 -29.000 ;
        RECT 216.680 -29.320 216.950 -29.050 ;
      LAYER met2 ;
        RECT 0.590 -29.410 217.040 -28.890 ;
    END
  END WL25
  PIN WL26
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER li1 ;
        RECT 7.340 -30.710 7.790 -30.260 ;
        RECT 20.840 -30.710 21.290 -30.260 ;
        RECT 34.340 -30.710 34.790 -30.260 ;
        RECT 47.840 -30.710 48.290 -30.260 ;
        RECT 61.340 -30.710 61.790 -30.260 ;
        RECT 74.840 -30.710 75.290 -30.260 ;
        RECT 88.340 -30.710 88.790 -30.260 ;
        RECT 101.840 -30.710 102.290 -30.260 ;
        RECT 115.340 -30.710 115.790 -30.260 ;
        RECT 128.840 -30.710 129.290 -30.260 ;
        RECT 142.340 -30.710 142.790 -30.260 ;
        RECT 155.840 -30.710 156.290 -30.260 ;
        RECT 169.340 -30.710 169.790 -30.260 ;
        RECT 182.840 -30.710 183.290 -30.260 ;
        RECT 196.340 -30.710 196.790 -30.260 ;
        RECT 209.840 -30.710 210.290 -30.260 ;
        RECT 0.590 -31.620 1.040 -31.180 ;
        RECT 14.090 -31.620 14.540 -31.180 ;
        RECT 27.590 -31.620 28.040 -31.180 ;
        RECT 41.090 -31.620 41.540 -31.180 ;
        RECT 54.590 -31.620 55.040 -31.180 ;
        RECT 68.090 -31.620 68.540 -31.180 ;
        RECT 81.590 -31.620 82.040 -31.180 ;
        RECT 95.090 -31.620 95.540 -31.180 ;
        RECT 108.590 -31.620 109.040 -31.180 ;
        RECT 122.090 -31.620 122.540 -31.180 ;
        RECT 135.590 -31.620 136.040 -31.180 ;
        RECT 149.090 -31.620 149.540 -31.180 ;
        RECT 162.590 -31.620 163.040 -31.180 ;
        RECT 176.090 -31.620 176.540 -31.180 ;
        RECT 189.590 -31.620 190.040 -31.180 ;
        RECT 203.090 -31.620 203.540 -31.180 ;
        RECT 216.590 -31.620 217.040 -31.180 ;
      LAYER mcon ;
        RECT 7.440 -30.610 7.690 -30.360 ;
        RECT 20.940 -30.610 21.190 -30.360 ;
        RECT 34.440 -30.610 34.690 -30.360 ;
        RECT 47.940 -30.610 48.190 -30.360 ;
        RECT 61.440 -30.610 61.690 -30.360 ;
        RECT 74.940 -30.610 75.190 -30.360 ;
        RECT 88.440 -30.610 88.690 -30.360 ;
        RECT 101.940 -30.610 102.190 -30.360 ;
        RECT 115.440 -30.610 115.690 -30.360 ;
        RECT 128.940 -30.610 129.190 -30.360 ;
        RECT 142.440 -30.610 142.690 -30.360 ;
        RECT 155.940 -30.610 156.190 -30.360 ;
        RECT 169.440 -30.610 169.690 -30.360 ;
        RECT 182.940 -30.610 183.190 -30.360 ;
        RECT 196.440 -30.610 196.690 -30.360 ;
        RECT 209.940 -30.610 210.190 -30.360 ;
        RECT 0.680 -31.530 0.950 -31.260 ;
        RECT 14.180 -31.530 14.450 -31.260 ;
        RECT 27.680 -31.530 27.950 -31.260 ;
        RECT 41.180 -31.530 41.450 -31.260 ;
        RECT 54.680 -31.530 54.950 -31.260 ;
        RECT 68.180 -31.530 68.450 -31.260 ;
        RECT 81.680 -31.530 81.950 -31.260 ;
        RECT 95.180 -31.530 95.450 -31.260 ;
        RECT 108.680 -31.530 108.950 -31.260 ;
        RECT 122.180 -31.530 122.450 -31.260 ;
        RECT 135.680 -31.530 135.950 -31.260 ;
        RECT 149.180 -31.530 149.450 -31.260 ;
        RECT 162.680 -31.530 162.950 -31.260 ;
        RECT 176.180 -31.530 176.450 -31.260 ;
        RECT 189.680 -31.530 189.950 -31.260 ;
        RECT 203.180 -31.530 203.450 -31.260 ;
        RECT 216.680 -31.530 216.950 -31.260 ;
      LAYER met1 ;
        RECT 0.590 -31.170 1.050 -30.700 ;
        RECT 0.580 -31.180 1.050 -31.170 ;
        RECT 7.330 -31.180 7.800 -30.250 ;
        RECT 0.580 -31.620 1.040 -31.180 ;
        RECT 14.080 -31.620 14.550 -30.700 ;
        RECT 20.830 -31.180 21.300 -30.250 ;
        RECT 27.580 -31.620 28.050 -30.700 ;
        RECT 34.330 -31.180 34.800 -30.250 ;
        RECT 41.080 -31.620 41.550 -30.700 ;
        RECT 47.830 -31.180 48.300 -30.250 ;
        RECT 54.580 -31.620 55.050 -30.700 ;
        RECT 61.330 -31.180 61.800 -30.250 ;
        RECT 68.080 -31.620 68.550 -30.700 ;
        RECT 74.830 -31.180 75.300 -30.250 ;
        RECT 81.580 -31.620 82.050 -30.700 ;
        RECT 88.330 -31.180 88.800 -30.250 ;
        RECT 95.080 -31.620 95.550 -30.700 ;
        RECT 101.830 -31.180 102.300 -30.250 ;
        RECT 108.580 -31.620 109.050 -30.700 ;
        RECT 115.330 -31.180 115.800 -30.250 ;
        RECT 122.080 -31.620 122.550 -30.700 ;
        RECT 128.830 -31.180 129.300 -30.250 ;
        RECT 135.580 -31.620 136.050 -30.700 ;
        RECT 142.330 -31.180 142.800 -30.250 ;
        RECT 149.080 -31.620 149.550 -30.700 ;
        RECT 155.830 -31.180 156.300 -30.250 ;
        RECT 162.580 -31.620 163.050 -30.700 ;
        RECT 169.330 -31.180 169.800 -30.250 ;
        RECT 176.080 -31.620 176.550 -30.700 ;
        RECT 182.830 -31.180 183.300 -30.250 ;
        RECT 189.580 -31.620 190.050 -30.700 ;
        RECT 196.330 -31.180 196.800 -30.250 ;
        RECT 203.080 -31.620 203.550 -30.700 ;
        RECT 209.830 -31.180 210.300 -30.250 ;
        RECT 216.580 -31.170 217.040 -30.700 ;
        RECT 216.580 -31.180 217.050 -31.170 ;
        RECT 216.590 -31.620 217.050 -31.180 ;
      LAYER via ;
        RECT 0.680 -31.030 0.950 -30.760 ;
        RECT 7.430 -31.050 7.700 -30.780 ;
        RECT 14.180 -31.030 14.450 -30.760 ;
        RECT 20.930 -31.080 21.200 -30.810 ;
        RECT 27.680 -31.030 27.950 -30.760 ;
        RECT 34.430 -31.080 34.700 -30.810 ;
        RECT 41.180 -31.030 41.450 -30.760 ;
        RECT 47.930 -31.050 48.200 -30.780 ;
        RECT 54.680 -31.030 54.950 -30.760 ;
        RECT 61.430 -31.050 61.700 -30.780 ;
        RECT 68.180 -31.030 68.450 -30.760 ;
        RECT 74.930 -31.080 75.200 -30.810 ;
        RECT 81.680 -31.030 81.950 -30.760 ;
        RECT 88.430 -31.080 88.700 -30.810 ;
        RECT 95.180 -31.030 95.450 -30.760 ;
        RECT 101.930 -31.050 102.200 -30.780 ;
        RECT 108.680 -31.030 108.950 -30.760 ;
        RECT 115.430 -31.050 115.700 -30.780 ;
        RECT 122.180 -31.030 122.450 -30.760 ;
        RECT 128.930 -31.080 129.200 -30.810 ;
        RECT 135.680 -31.030 135.950 -30.760 ;
        RECT 142.430 -31.080 142.700 -30.810 ;
        RECT 149.180 -31.030 149.450 -30.760 ;
        RECT 155.930 -31.050 156.200 -30.780 ;
        RECT 162.680 -31.030 162.950 -30.760 ;
        RECT 169.430 -31.050 169.700 -30.780 ;
        RECT 176.180 -31.030 176.450 -30.760 ;
        RECT 182.930 -31.080 183.200 -30.810 ;
        RECT 189.680 -31.030 189.950 -30.760 ;
        RECT 196.430 -31.080 196.700 -30.810 ;
        RECT 203.180 -31.030 203.450 -30.760 ;
        RECT 209.930 -31.050 210.200 -30.780 ;
        RECT 216.680 -31.030 216.950 -30.760 ;
      LAYER met2 ;
        RECT 0.580 -30.660 1.060 -30.650 ;
        RECT 108.570 -30.660 109.060 -30.650 ;
        RECT 216.570 -30.660 217.050 -30.650 ;
        RECT 0.580 -30.670 14.590 -30.660 ;
        RECT 41.040 -30.670 68.590 -30.660 ;
        RECT 95.040 -30.670 122.590 -30.660 ;
        RECT 149.040 -30.670 176.590 -30.660 ;
        RECT 203.040 -30.670 217.050 -30.660 ;
        RECT 0.580 -31.170 217.050 -30.670 ;
        RECT 0.590 -31.180 217.040 -31.170 ;
        RECT 14.040 -31.190 41.590 -31.180 ;
        RECT 68.040 -31.190 95.590 -31.180 ;
        RECT 122.040 -31.190 149.590 -31.180 ;
        RECT 176.040 -31.190 203.590 -31.180 ;
    END
  END WL26
  PIN WL27
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER li1 ;
        RECT 0.590 -32.510 1.040 -32.070 ;
        RECT 14.090 -32.510 14.540 -32.070 ;
        RECT 27.590 -32.510 28.040 -32.070 ;
        RECT 41.090 -32.510 41.540 -32.070 ;
        RECT 54.590 -32.510 55.040 -32.070 ;
        RECT 68.090 -32.510 68.540 -32.070 ;
        RECT 81.590 -32.510 82.040 -32.070 ;
        RECT 95.090 -32.510 95.540 -32.070 ;
        RECT 108.590 -32.510 109.040 -32.070 ;
        RECT 122.090 -32.510 122.540 -32.070 ;
        RECT 135.590 -32.510 136.040 -32.070 ;
        RECT 149.090 -32.510 149.540 -32.070 ;
        RECT 162.590 -32.510 163.040 -32.070 ;
        RECT 176.090 -32.510 176.540 -32.070 ;
        RECT 189.590 -32.510 190.040 -32.070 ;
        RECT 203.090 -32.510 203.540 -32.070 ;
        RECT 216.590 -32.510 217.040 -32.070 ;
        RECT 7.340 -33.430 7.790 -32.980 ;
        RECT 20.840 -33.430 21.290 -32.980 ;
        RECT 34.340 -33.430 34.790 -32.980 ;
        RECT 47.840 -33.430 48.290 -32.980 ;
        RECT 61.340 -33.430 61.790 -32.980 ;
        RECT 74.840 -33.430 75.290 -32.980 ;
        RECT 88.340 -33.430 88.790 -32.980 ;
        RECT 101.840 -33.430 102.290 -32.980 ;
        RECT 115.340 -33.430 115.790 -32.980 ;
        RECT 128.840 -33.430 129.290 -32.980 ;
        RECT 142.340 -33.430 142.790 -32.980 ;
        RECT 155.840 -33.430 156.290 -32.980 ;
        RECT 169.340 -33.430 169.790 -32.980 ;
        RECT 182.840 -33.430 183.290 -32.980 ;
        RECT 196.340 -33.430 196.790 -32.980 ;
        RECT 209.840 -33.430 210.290 -32.980 ;
      LAYER mcon ;
        RECT 0.680 -32.430 0.950 -32.160 ;
        RECT 14.180 -32.430 14.450 -32.160 ;
        RECT 27.680 -32.430 27.950 -32.160 ;
        RECT 41.180 -32.430 41.450 -32.160 ;
        RECT 54.680 -32.430 54.950 -32.160 ;
        RECT 68.180 -32.430 68.450 -32.160 ;
        RECT 81.680 -32.430 81.950 -32.160 ;
        RECT 95.180 -32.430 95.450 -32.160 ;
        RECT 108.680 -32.430 108.950 -32.160 ;
        RECT 122.180 -32.430 122.450 -32.160 ;
        RECT 135.680 -32.430 135.950 -32.160 ;
        RECT 149.180 -32.430 149.450 -32.160 ;
        RECT 162.680 -32.430 162.950 -32.160 ;
        RECT 176.180 -32.430 176.450 -32.160 ;
        RECT 189.680 -32.430 189.950 -32.160 ;
        RECT 203.180 -32.430 203.450 -32.160 ;
        RECT 216.680 -32.430 216.950 -32.160 ;
        RECT 7.440 -33.330 7.690 -33.080 ;
        RECT 20.940 -33.330 21.190 -33.080 ;
        RECT 34.440 -33.330 34.690 -33.080 ;
        RECT 47.940 -33.330 48.190 -33.080 ;
        RECT 61.440 -33.330 61.690 -33.080 ;
        RECT 74.940 -33.330 75.190 -33.080 ;
        RECT 88.440 -33.330 88.690 -33.080 ;
        RECT 101.940 -33.330 102.190 -33.080 ;
        RECT 115.440 -33.330 115.690 -33.080 ;
        RECT 128.940 -33.330 129.190 -33.080 ;
        RECT 142.440 -33.330 142.690 -33.080 ;
        RECT 155.940 -33.330 156.190 -33.080 ;
        RECT 169.440 -33.330 169.690 -33.080 ;
        RECT 182.940 -33.330 183.190 -33.080 ;
        RECT 196.440 -33.330 196.690 -33.080 ;
        RECT 209.940 -33.330 210.190 -33.080 ;
      LAYER met1 ;
        RECT 0.580 -32.510 1.040 -32.070 ;
        RECT 0.580 -32.520 1.050 -32.510 ;
        RECT 0.590 -32.990 1.050 -32.520 ;
        RECT 7.330 -33.440 7.800 -32.510 ;
        RECT 14.080 -32.990 14.550 -32.070 ;
        RECT 20.830 -33.440 21.300 -32.510 ;
        RECT 27.580 -32.990 28.050 -32.070 ;
        RECT 34.330 -33.440 34.800 -32.510 ;
        RECT 41.080 -32.990 41.550 -32.070 ;
        RECT 47.830 -33.440 48.300 -32.510 ;
        RECT 54.580 -32.990 55.050 -32.070 ;
        RECT 61.330 -33.440 61.800 -32.510 ;
        RECT 68.080 -32.990 68.550 -32.070 ;
        RECT 74.830 -33.440 75.300 -32.510 ;
        RECT 81.580 -32.990 82.050 -32.070 ;
        RECT 88.330 -33.440 88.800 -32.510 ;
        RECT 95.080 -32.990 95.550 -32.070 ;
        RECT 101.830 -33.440 102.300 -32.510 ;
        RECT 108.580 -32.990 109.050 -32.070 ;
        RECT 115.330 -33.440 115.800 -32.510 ;
        RECT 122.080 -32.990 122.550 -32.070 ;
        RECT 128.830 -33.440 129.300 -32.510 ;
        RECT 135.580 -32.990 136.050 -32.070 ;
        RECT 142.330 -33.440 142.800 -32.510 ;
        RECT 149.080 -32.990 149.550 -32.070 ;
        RECT 155.830 -33.440 156.300 -32.510 ;
        RECT 162.580 -32.990 163.050 -32.070 ;
        RECT 169.330 -33.440 169.800 -32.510 ;
        RECT 176.080 -32.990 176.550 -32.070 ;
        RECT 182.830 -33.440 183.300 -32.510 ;
        RECT 189.580 -32.990 190.050 -32.070 ;
        RECT 196.330 -33.440 196.800 -32.510 ;
        RECT 203.080 -32.990 203.550 -32.070 ;
        RECT 216.590 -32.510 217.050 -32.070 ;
        RECT 209.830 -33.440 210.300 -32.510 ;
        RECT 216.580 -32.520 217.050 -32.510 ;
        RECT 216.580 -32.990 217.040 -32.520 ;
      LAYER via ;
        RECT 0.680 -32.930 0.950 -32.660 ;
        RECT 7.430 -32.880 7.700 -32.610 ;
        RECT 14.180 -32.930 14.450 -32.660 ;
        RECT 20.930 -32.910 21.200 -32.640 ;
        RECT 27.680 -32.930 27.950 -32.660 ;
        RECT 34.430 -32.910 34.700 -32.640 ;
        RECT 41.180 -32.930 41.450 -32.660 ;
        RECT 47.930 -32.880 48.200 -32.610 ;
        RECT 54.680 -32.930 54.950 -32.660 ;
        RECT 61.430 -32.880 61.700 -32.610 ;
        RECT 68.180 -32.930 68.450 -32.660 ;
        RECT 74.930 -32.910 75.200 -32.640 ;
        RECT 81.680 -32.930 81.950 -32.660 ;
        RECT 88.430 -32.910 88.700 -32.640 ;
        RECT 95.180 -32.930 95.450 -32.660 ;
        RECT 101.930 -32.880 102.200 -32.610 ;
        RECT 108.680 -32.930 108.950 -32.660 ;
        RECT 115.430 -32.880 115.700 -32.610 ;
        RECT 122.180 -32.930 122.450 -32.660 ;
        RECT 128.930 -32.910 129.200 -32.640 ;
        RECT 135.680 -32.930 135.950 -32.660 ;
        RECT 142.430 -32.910 142.700 -32.640 ;
        RECT 149.180 -32.930 149.450 -32.660 ;
        RECT 155.930 -32.880 156.200 -32.610 ;
        RECT 162.680 -32.930 162.950 -32.660 ;
        RECT 169.430 -32.880 169.700 -32.610 ;
        RECT 176.180 -32.930 176.450 -32.660 ;
        RECT 182.930 -32.910 183.200 -32.640 ;
        RECT 189.680 -32.930 189.950 -32.660 ;
        RECT 196.430 -32.910 196.700 -32.640 ;
        RECT 203.180 -32.930 203.450 -32.660 ;
        RECT 209.930 -32.880 210.200 -32.610 ;
        RECT 216.680 -32.930 216.950 -32.660 ;
      LAYER met2 ;
        RECT 0.590 -32.510 14.590 -32.500 ;
        RECT 41.040 -32.510 68.590 -32.500 ;
        RECT 95.040 -32.510 122.590 -32.500 ;
        RECT 149.040 -32.510 176.590 -32.500 ;
        RECT 203.040 -32.510 217.040 -32.500 ;
        RECT 0.590 -32.520 217.040 -32.510 ;
        RECT 0.580 -33.020 217.050 -32.520 ;
        RECT 0.580 -33.030 1.060 -33.020 ;
        RECT 14.040 -33.030 41.590 -33.020 ;
        RECT 68.040 -33.030 95.590 -33.020 ;
        RECT 108.570 -33.030 109.060 -33.020 ;
        RECT 122.040 -33.030 149.590 -33.020 ;
        RECT 176.040 -33.030 203.590 -33.020 ;
        RECT 216.570 -33.030 217.050 -33.020 ;
    END
  END WL27
  PIN WL28
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER li1 ;
        RECT 7.340 -34.320 7.790 -33.870 ;
        RECT 20.840 -34.320 21.290 -33.870 ;
        RECT 34.340 -34.320 34.790 -33.870 ;
        RECT 47.840 -34.320 48.290 -33.870 ;
        RECT 61.340 -34.320 61.790 -33.870 ;
        RECT 74.840 -34.320 75.290 -33.870 ;
        RECT 88.340 -34.320 88.790 -33.870 ;
        RECT 101.840 -34.320 102.290 -33.870 ;
        RECT 115.340 -34.320 115.790 -33.870 ;
        RECT 128.840 -34.320 129.290 -33.870 ;
        RECT 142.340 -34.320 142.790 -33.870 ;
        RECT 155.840 -34.320 156.290 -33.870 ;
        RECT 169.340 -34.320 169.790 -33.870 ;
        RECT 182.840 -34.320 183.290 -33.870 ;
        RECT 196.340 -34.320 196.790 -33.870 ;
        RECT 209.840 -34.320 210.290 -33.870 ;
        RECT 0.590 -35.230 1.040 -34.790 ;
        RECT 14.090 -35.230 14.540 -34.790 ;
        RECT 27.590 -35.230 28.040 -34.790 ;
        RECT 41.090 -35.230 41.540 -34.790 ;
        RECT 54.590 -35.230 55.040 -34.790 ;
        RECT 68.090 -35.230 68.540 -34.790 ;
        RECT 81.590 -35.230 82.040 -34.790 ;
        RECT 95.090 -35.230 95.540 -34.790 ;
        RECT 108.590 -35.230 109.040 -34.790 ;
        RECT 122.090 -35.230 122.540 -34.790 ;
        RECT 135.590 -35.230 136.040 -34.790 ;
        RECT 149.090 -35.230 149.540 -34.790 ;
        RECT 162.590 -35.230 163.040 -34.790 ;
        RECT 176.090 -35.230 176.540 -34.790 ;
        RECT 189.590 -35.230 190.040 -34.790 ;
        RECT 203.090 -35.230 203.540 -34.790 ;
        RECT 216.590 -35.230 217.040 -34.790 ;
      LAYER mcon ;
        RECT 7.440 -34.220 7.690 -33.970 ;
        RECT 20.940 -34.220 21.190 -33.970 ;
        RECT 34.440 -34.220 34.690 -33.970 ;
        RECT 47.940 -34.220 48.190 -33.970 ;
        RECT 61.440 -34.220 61.690 -33.970 ;
        RECT 74.940 -34.220 75.190 -33.970 ;
        RECT 88.440 -34.220 88.690 -33.970 ;
        RECT 101.940 -34.220 102.190 -33.970 ;
        RECT 115.440 -34.220 115.690 -33.970 ;
        RECT 128.940 -34.220 129.190 -33.970 ;
        RECT 142.440 -34.220 142.690 -33.970 ;
        RECT 155.940 -34.220 156.190 -33.970 ;
        RECT 169.440 -34.220 169.690 -33.970 ;
        RECT 182.940 -34.220 183.190 -33.970 ;
        RECT 196.440 -34.220 196.690 -33.970 ;
        RECT 209.940 -34.220 210.190 -33.970 ;
        RECT 0.680 -35.140 0.950 -34.870 ;
        RECT 14.180 -35.140 14.450 -34.870 ;
        RECT 27.680 -35.140 27.950 -34.870 ;
        RECT 41.180 -35.140 41.450 -34.870 ;
        RECT 54.680 -35.140 54.950 -34.870 ;
        RECT 68.180 -35.140 68.450 -34.870 ;
        RECT 81.680 -35.140 81.950 -34.870 ;
        RECT 95.180 -35.140 95.450 -34.870 ;
        RECT 108.680 -35.140 108.950 -34.870 ;
        RECT 122.180 -35.140 122.450 -34.870 ;
        RECT 135.680 -35.140 135.950 -34.870 ;
        RECT 149.180 -35.140 149.450 -34.870 ;
        RECT 162.680 -35.140 162.950 -34.870 ;
        RECT 176.180 -35.140 176.450 -34.870 ;
        RECT 189.680 -35.140 189.950 -34.870 ;
        RECT 203.180 -35.140 203.450 -34.870 ;
        RECT 216.680 -35.140 216.950 -34.870 ;
      LAYER met1 ;
        RECT 0.590 -34.780 1.050 -34.310 ;
        RECT 0.580 -34.790 1.050 -34.780 ;
        RECT 7.330 -34.790 7.800 -33.860 ;
        RECT 0.580 -35.230 1.040 -34.790 ;
        RECT 14.080 -35.230 14.550 -34.310 ;
        RECT 20.830 -34.790 21.300 -33.860 ;
        RECT 27.580 -35.230 28.050 -34.310 ;
        RECT 34.330 -34.790 34.800 -33.860 ;
        RECT 41.080 -35.230 41.550 -34.310 ;
        RECT 47.830 -34.790 48.300 -33.860 ;
        RECT 54.580 -35.230 55.050 -34.310 ;
        RECT 61.330 -34.790 61.800 -33.860 ;
        RECT 68.080 -35.230 68.550 -34.310 ;
        RECT 74.830 -34.790 75.300 -33.860 ;
        RECT 81.580 -35.230 82.050 -34.310 ;
        RECT 88.330 -34.790 88.800 -33.860 ;
        RECT 95.080 -35.230 95.550 -34.310 ;
        RECT 101.830 -34.790 102.300 -33.860 ;
        RECT 108.580 -35.230 109.050 -34.310 ;
        RECT 115.330 -34.790 115.800 -33.860 ;
        RECT 122.080 -35.230 122.550 -34.310 ;
        RECT 128.830 -34.790 129.300 -33.860 ;
        RECT 135.580 -35.230 136.050 -34.310 ;
        RECT 142.330 -34.790 142.800 -33.860 ;
        RECT 149.080 -35.230 149.550 -34.310 ;
        RECT 155.830 -34.790 156.300 -33.860 ;
        RECT 162.580 -35.230 163.050 -34.310 ;
        RECT 169.330 -34.790 169.800 -33.860 ;
        RECT 176.080 -35.230 176.550 -34.310 ;
        RECT 182.830 -34.790 183.300 -33.860 ;
        RECT 189.580 -35.230 190.050 -34.310 ;
        RECT 196.330 -34.790 196.800 -33.860 ;
        RECT 203.080 -35.230 203.550 -34.310 ;
        RECT 209.830 -34.790 210.300 -33.860 ;
        RECT 216.580 -34.780 217.040 -34.310 ;
        RECT 216.580 -34.790 217.050 -34.780 ;
        RECT 216.590 -35.230 217.050 -34.790 ;
      LAYER via ;
        RECT 0.680 -34.640 0.950 -34.370 ;
        RECT 7.430 -34.690 7.700 -34.420 ;
        RECT 14.180 -34.640 14.450 -34.370 ;
        RECT 20.930 -34.660 21.200 -34.390 ;
        RECT 27.680 -34.640 27.950 -34.370 ;
        RECT 34.430 -34.660 34.700 -34.390 ;
        RECT 41.180 -34.640 41.450 -34.370 ;
        RECT 47.930 -34.690 48.200 -34.420 ;
        RECT 54.680 -34.640 54.950 -34.370 ;
        RECT 61.430 -34.690 61.700 -34.420 ;
        RECT 68.180 -34.640 68.450 -34.370 ;
        RECT 74.930 -34.660 75.200 -34.390 ;
        RECT 81.680 -34.640 81.950 -34.370 ;
        RECT 88.430 -34.660 88.700 -34.390 ;
        RECT 95.180 -34.640 95.450 -34.370 ;
        RECT 101.930 -34.690 102.200 -34.420 ;
        RECT 108.680 -34.640 108.950 -34.370 ;
        RECT 115.430 -34.690 115.700 -34.420 ;
        RECT 122.180 -34.640 122.450 -34.370 ;
        RECT 128.930 -34.660 129.200 -34.390 ;
        RECT 135.680 -34.640 135.950 -34.370 ;
        RECT 142.430 -34.660 142.700 -34.390 ;
        RECT 149.180 -34.640 149.450 -34.370 ;
        RECT 155.930 -34.690 156.200 -34.420 ;
        RECT 162.680 -34.640 162.950 -34.370 ;
        RECT 169.430 -34.690 169.700 -34.420 ;
        RECT 176.180 -34.640 176.450 -34.370 ;
        RECT 182.930 -34.660 183.200 -34.390 ;
        RECT 189.680 -34.640 189.950 -34.370 ;
        RECT 196.430 -34.660 196.700 -34.390 ;
        RECT 203.180 -34.640 203.450 -34.370 ;
        RECT 209.930 -34.690 210.200 -34.420 ;
        RECT 216.680 -34.640 216.950 -34.370 ;
      LAYER met2 ;
        RECT 14.040 -34.280 41.590 -34.270 ;
        RECT 68.040 -34.280 95.590 -34.270 ;
        RECT 122.040 -34.280 149.590 -34.270 ;
        RECT 176.040 -34.280 203.590 -34.270 ;
        RECT 0.590 -34.290 217.040 -34.280 ;
        RECT 0.580 -34.770 217.050 -34.290 ;
        RECT 0.590 -34.790 217.040 -34.770 ;
        RECT 0.590 -34.800 14.590 -34.790 ;
        RECT 41.040 -34.800 68.590 -34.790 ;
        RECT 95.040 -34.800 122.590 -34.790 ;
        RECT 149.040 -34.800 176.590 -34.790 ;
        RECT 203.040 -34.800 217.040 -34.790 ;
    END
  END WL28
  PIN WL29
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER li1 ;
        RECT 0.590 -36.120 1.040 -35.680 ;
        RECT 14.090 -36.120 14.540 -35.680 ;
        RECT 27.590 -36.120 28.040 -35.680 ;
        RECT 41.090 -36.120 41.540 -35.680 ;
        RECT 54.590 -36.120 55.040 -35.680 ;
        RECT 68.090 -36.120 68.540 -35.680 ;
        RECT 81.590 -36.120 82.040 -35.680 ;
        RECT 95.090 -36.120 95.540 -35.680 ;
        RECT 108.590 -36.120 109.040 -35.680 ;
        RECT 122.090 -36.120 122.540 -35.680 ;
        RECT 135.590 -36.120 136.040 -35.680 ;
        RECT 149.090 -36.120 149.540 -35.680 ;
        RECT 162.590 -36.120 163.040 -35.680 ;
        RECT 176.090 -36.120 176.540 -35.680 ;
        RECT 189.590 -36.120 190.040 -35.680 ;
        RECT 203.090 -36.120 203.540 -35.680 ;
        RECT 216.590 -36.120 217.040 -35.680 ;
        RECT 7.340 -37.040 7.790 -36.590 ;
        RECT 20.840 -37.040 21.290 -36.590 ;
        RECT 34.340 -37.040 34.790 -36.590 ;
        RECT 47.840 -37.040 48.290 -36.590 ;
        RECT 61.340 -37.040 61.790 -36.590 ;
        RECT 74.840 -37.040 75.290 -36.590 ;
        RECT 88.340 -37.040 88.790 -36.590 ;
        RECT 101.840 -37.040 102.290 -36.590 ;
        RECT 115.340 -37.040 115.790 -36.590 ;
        RECT 128.840 -37.040 129.290 -36.590 ;
        RECT 142.340 -37.040 142.790 -36.590 ;
        RECT 155.840 -37.040 156.290 -36.590 ;
        RECT 169.340 -37.040 169.790 -36.590 ;
        RECT 182.840 -37.040 183.290 -36.590 ;
        RECT 196.340 -37.040 196.790 -36.590 ;
        RECT 209.840 -37.040 210.290 -36.590 ;
      LAYER mcon ;
        RECT 0.680 -36.040 0.950 -35.770 ;
        RECT 14.180 -36.040 14.450 -35.770 ;
        RECT 27.680 -36.040 27.950 -35.770 ;
        RECT 41.180 -36.040 41.450 -35.770 ;
        RECT 54.680 -36.040 54.950 -35.770 ;
        RECT 68.180 -36.040 68.450 -35.770 ;
        RECT 81.680 -36.040 81.950 -35.770 ;
        RECT 95.180 -36.040 95.450 -35.770 ;
        RECT 108.680 -36.040 108.950 -35.770 ;
        RECT 122.180 -36.040 122.450 -35.770 ;
        RECT 135.680 -36.040 135.950 -35.770 ;
        RECT 149.180 -36.040 149.450 -35.770 ;
        RECT 162.680 -36.040 162.950 -35.770 ;
        RECT 176.180 -36.040 176.450 -35.770 ;
        RECT 189.680 -36.040 189.950 -35.770 ;
        RECT 203.180 -36.040 203.450 -35.770 ;
        RECT 216.680 -36.040 216.950 -35.770 ;
        RECT 7.440 -36.940 7.690 -36.690 ;
        RECT 20.940 -36.940 21.190 -36.690 ;
        RECT 34.440 -36.940 34.690 -36.690 ;
        RECT 47.940 -36.940 48.190 -36.690 ;
        RECT 61.440 -36.940 61.690 -36.690 ;
        RECT 74.940 -36.940 75.190 -36.690 ;
        RECT 88.440 -36.940 88.690 -36.690 ;
        RECT 101.940 -36.940 102.190 -36.690 ;
        RECT 115.440 -36.940 115.690 -36.690 ;
        RECT 128.940 -36.940 129.190 -36.690 ;
        RECT 142.440 -36.940 142.690 -36.690 ;
        RECT 155.940 -36.940 156.190 -36.690 ;
        RECT 169.440 -36.940 169.690 -36.690 ;
        RECT 182.940 -36.940 183.190 -36.690 ;
        RECT 196.440 -36.940 196.690 -36.690 ;
        RECT 209.940 -36.940 210.190 -36.690 ;
      LAYER met1 ;
        RECT 0.580 -36.120 1.040 -35.680 ;
        RECT 0.580 -36.130 1.050 -36.120 ;
        RECT 0.590 -36.600 1.050 -36.130 ;
        RECT 7.330 -37.050 7.800 -36.120 ;
        RECT 14.080 -36.600 14.550 -35.680 ;
        RECT 20.830 -37.050 21.300 -36.120 ;
        RECT 27.580 -36.600 28.050 -35.680 ;
        RECT 34.330 -37.050 34.800 -36.120 ;
        RECT 41.080 -36.600 41.550 -35.680 ;
        RECT 47.830 -37.050 48.300 -36.120 ;
        RECT 54.580 -36.600 55.050 -35.680 ;
        RECT 61.330 -37.050 61.800 -36.120 ;
        RECT 68.080 -36.600 68.550 -35.680 ;
        RECT 74.830 -37.050 75.300 -36.120 ;
        RECT 81.580 -36.600 82.050 -35.680 ;
        RECT 88.330 -37.050 88.800 -36.120 ;
        RECT 95.080 -36.600 95.550 -35.680 ;
        RECT 101.830 -37.050 102.300 -36.120 ;
        RECT 108.580 -36.600 109.050 -35.680 ;
        RECT 115.330 -37.050 115.800 -36.120 ;
        RECT 122.080 -36.600 122.550 -35.680 ;
        RECT 128.830 -37.050 129.300 -36.120 ;
        RECT 135.580 -36.600 136.050 -35.680 ;
        RECT 142.330 -37.050 142.800 -36.120 ;
        RECT 149.080 -36.600 149.550 -35.680 ;
        RECT 155.830 -37.050 156.300 -36.120 ;
        RECT 162.580 -36.600 163.050 -35.680 ;
        RECT 169.330 -37.050 169.800 -36.120 ;
        RECT 176.080 -36.600 176.550 -35.680 ;
        RECT 182.830 -37.050 183.300 -36.120 ;
        RECT 189.580 -36.600 190.050 -35.680 ;
        RECT 196.330 -37.050 196.800 -36.120 ;
        RECT 203.080 -36.600 203.550 -35.680 ;
        RECT 216.590 -36.120 217.050 -35.680 ;
        RECT 209.830 -37.050 210.300 -36.120 ;
        RECT 216.580 -36.130 217.050 -36.120 ;
        RECT 216.580 -36.600 217.040 -36.130 ;
      LAYER via ;
        RECT 0.680 -36.540 0.950 -36.270 ;
        RECT 7.430 -36.520 7.700 -36.250 ;
        RECT 14.180 -36.540 14.450 -36.270 ;
        RECT 20.930 -36.490 21.200 -36.220 ;
        RECT 27.680 -36.540 27.950 -36.270 ;
        RECT 34.430 -36.490 34.700 -36.220 ;
        RECT 41.180 -36.540 41.450 -36.270 ;
        RECT 47.930 -36.520 48.200 -36.250 ;
        RECT 54.680 -36.540 54.950 -36.270 ;
        RECT 61.430 -36.520 61.700 -36.250 ;
        RECT 68.180 -36.540 68.450 -36.270 ;
        RECT 74.930 -36.490 75.200 -36.220 ;
        RECT 81.680 -36.540 81.950 -36.270 ;
        RECT 88.430 -36.490 88.700 -36.220 ;
        RECT 95.180 -36.540 95.450 -36.270 ;
        RECT 101.930 -36.520 102.200 -36.250 ;
        RECT 108.680 -36.540 108.950 -36.270 ;
        RECT 115.430 -36.520 115.700 -36.250 ;
        RECT 122.180 -36.540 122.450 -36.270 ;
        RECT 128.930 -36.490 129.200 -36.220 ;
        RECT 135.680 -36.540 135.950 -36.270 ;
        RECT 142.430 -36.490 142.700 -36.220 ;
        RECT 149.180 -36.540 149.450 -36.270 ;
        RECT 155.930 -36.520 156.200 -36.250 ;
        RECT 162.680 -36.540 162.950 -36.270 ;
        RECT 169.430 -36.520 169.700 -36.250 ;
        RECT 176.180 -36.540 176.450 -36.270 ;
        RECT 182.930 -36.490 183.200 -36.220 ;
        RECT 189.680 -36.540 189.950 -36.270 ;
        RECT 196.430 -36.490 196.700 -36.220 ;
        RECT 203.180 -36.540 203.450 -36.270 ;
        RECT 209.930 -36.520 210.200 -36.250 ;
        RECT 216.680 -36.540 216.950 -36.270 ;
      LAYER met2 ;
        RECT 14.040 -36.120 41.590 -36.110 ;
        RECT 68.040 -36.120 95.590 -36.110 ;
        RECT 122.040 -36.120 149.590 -36.110 ;
        RECT 176.040 -36.120 203.590 -36.110 ;
        RECT 0.590 -36.130 217.040 -36.120 ;
        RECT 0.580 -36.610 217.050 -36.130 ;
        RECT 0.590 -36.630 217.040 -36.610 ;
        RECT 0.590 -36.640 14.590 -36.630 ;
        RECT 41.040 -36.640 68.590 -36.630 ;
        RECT 95.040 -36.640 122.590 -36.630 ;
        RECT 149.040 -36.640 176.590 -36.630 ;
        RECT 203.040 -36.640 217.040 -36.630 ;
        RECT 0.590 -36.650 1.070 -36.640 ;
        RECT 108.560 -36.650 109.070 -36.640 ;
        RECT 216.560 -36.650 217.040 -36.640 ;
    END
  END WL29
  PIN WL30
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER li1 ;
        RECT 7.340 -37.930 7.790 -37.480 ;
        RECT 20.840 -37.930 21.290 -37.480 ;
        RECT 34.340 -37.930 34.790 -37.480 ;
        RECT 47.840 -37.930 48.290 -37.480 ;
        RECT 61.340 -37.930 61.790 -37.480 ;
        RECT 74.840 -37.930 75.290 -37.480 ;
        RECT 88.340 -37.930 88.790 -37.480 ;
        RECT 101.840 -37.930 102.290 -37.480 ;
        RECT 115.340 -37.930 115.790 -37.480 ;
        RECT 128.840 -37.930 129.290 -37.480 ;
        RECT 142.340 -37.930 142.790 -37.480 ;
        RECT 155.840 -37.930 156.290 -37.480 ;
        RECT 169.340 -37.930 169.790 -37.480 ;
        RECT 182.840 -37.930 183.290 -37.480 ;
        RECT 196.340 -37.930 196.790 -37.480 ;
        RECT 209.840 -37.930 210.290 -37.480 ;
        RECT 0.590 -38.840 1.040 -38.400 ;
        RECT 14.090 -38.840 14.540 -38.400 ;
        RECT 27.590 -38.840 28.040 -38.400 ;
        RECT 41.090 -38.840 41.540 -38.400 ;
        RECT 54.590 -38.840 55.040 -38.400 ;
        RECT 68.090 -38.840 68.540 -38.400 ;
        RECT 81.590 -38.840 82.040 -38.400 ;
        RECT 95.090 -38.840 95.540 -38.400 ;
        RECT 108.590 -38.840 109.040 -38.400 ;
        RECT 122.090 -38.840 122.540 -38.400 ;
        RECT 135.590 -38.840 136.040 -38.400 ;
        RECT 149.090 -38.840 149.540 -38.400 ;
        RECT 162.590 -38.840 163.040 -38.400 ;
        RECT 176.090 -38.840 176.540 -38.400 ;
        RECT 189.590 -38.840 190.040 -38.400 ;
        RECT 203.090 -38.840 203.540 -38.400 ;
        RECT 216.590 -38.840 217.040 -38.400 ;
      LAYER mcon ;
        RECT 7.440 -37.830 7.690 -37.580 ;
        RECT 20.940 -37.830 21.190 -37.580 ;
        RECT 34.440 -37.830 34.690 -37.580 ;
        RECT 47.940 -37.830 48.190 -37.580 ;
        RECT 61.440 -37.830 61.690 -37.580 ;
        RECT 74.940 -37.830 75.190 -37.580 ;
        RECT 88.440 -37.830 88.690 -37.580 ;
        RECT 101.940 -37.830 102.190 -37.580 ;
        RECT 115.440 -37.830 115.690 -37.580 ;
        RECT 128.940 -37.830 129.190 -37.580 ;
        RECT 142.440 -37.830 142.690 -37.580 ;
        RECT 155.940 -37.830 156.190 -37.580 ;
        RECT 169.440 -37.830 169.690 -37.580 ;
        RECT 182.940 -37.830 183.190 -37.580 ;
        RECT 196.440 -37.830 196.690 -37.580 ;
        RECT 209.940 -37.830 210.190 -37.580 ;
        RECT 0.680 -38.750 0.950 -38.480 ;
        RECT 14.180 -38.750 14.450 -38.480 ;
        RECT 27.680 -38.750 27.950 -38.480 ;
        RECT 41.180 -38.750 41.450 -38.480 ;
        RECT 54.680 -38.750 54.950 -38.480 ;
        RECT 68.180 -38.750 68.450 -38.480 ;
        RECT 81.680 -38.750 81.950 -38.480 ;
        RECT 95.180 -38.750 95.450 -38.480 ;
        RECT 108.680 -38.750 108.950 -38.480 ;
        RECT 122.180 -38.750 122.450 -38.480 ;
        RECT 135.680 -38.750 135.950 -38.480 ;
        RECT 149.180 -38.750 149.450 -38.480 ;
        RECT 162.680 -38.750 162.950 -38.480 ;
        RECT 176.180 -38.750 176.450 -38.480 ;
        RECT 189.680 -38.750 189.950 -38.480 ;
        RECT 203.180 -38.750 203.450 -38.480 ;
        RECT 216.680 -38.750 216.950 -38.480 ;
      LAYER met1 ;
        RECT 0.590 -38.390 1.050 -37.920 ;
        RECT 0.580 -38.400 1.050 -38.390 ;
        RECT 7.330 -38.400 7.800 -37.470 ;
        RECT 0.580 -38.840 1.040 -38.400 ;
        RECT 14.080 -38.840 14.550 -37.920 ;
        RECT 20.830 -38.400 21.300 -37.470 ;
        RECT 27.580 -38.840 28.050 -37.920 ;
        RECT 34.330 -38.400 34.800 -37.470 ;
        RECT 41.080 -38.840 41.550 -37.920 ;
        RECT 47.830 -38.400 48.300 -37.470 ;
        RECT 54.580 -38.840 55.050 -37.920 ;
        RECT 61.330 -38.400 61.800 -37.470 ;
        RECT 68.080 -38.840 68.550 -37.920 ;
        RECT 74.830 -38.400 75.300 -37.470 ;
        RECT 81.580 -38.840 82.050 -37.920 ;
        RECT 88.330 -38.400 88.800 -37.470 ;
        RECT 95.080 -38.840 95.550 -37.920 ;
        RECT 101.830 -38.400 102.300 -37.470 ;
        RECT 108.580 -38.840 109.050 -37.920 ;
        RECT 115.330 -38.400 115.800 -37.470 ;
        RECT 122.080 -38.840 122.550 -37.920 ;
        RECT 128.830 -38.400 129.300 -37.470 ;
        RECT 135.580 -38.840 136.050 -37.920 ;
        RECT 142.330 -38.400 142.800 -37.470 ;
        RECT 149.080 -38.840 149.550 -37.920 ;
        RECT 155.830 -38.400 156.300 -37.470 ;
        RECT 162.580 -38.840 163.050 -37.920 ;
        RECT 169.330 -38.400 169.800 -37.470 ;
        RECT 176.080 -38.840 176.550 -37.920 ;
        RECT 182.830 -38.400 183.300 -37.470 ;
        RECT 189.580 -38.840 190.050 -37.920 ;
        RECT 196.330 -38.400 196.800 -37.470 ;
        RECT 203.080 -38.840 203.550 -37.920 ;
        RECT 209.830 -38.400 210.300 -37.470 ;
        RECT 216.580 -38.390 217.040 -37.920 ;
        RECT 216.580 -38.400 217.050 -38.390 ;
        RECT 216.590 -38.840 217.050 -38.400 ;
      LAYER via ;
        RECT 0.680 -38.250 0.950 -37.980 ;
        RECT 7.430 -38.300 7.700 -38.030 ;
        RECT 14.180 -38.250 14.450 -37.980 ;
        RECT 20.930 -38.300 21.200 -38.030 ;
        RECT 27.680 -38.250 27.950 -37.980 ;
        RECT 34.430 -38.300 34.700 -38.030 ;
        RECT 41.180 -38.250 41.450 -37.980 ;
        RECT 47.930 -38.300 48.200 -38.030 ;
        RECT 54.680 -38.250 54.950 -37.980 ;
        RECT 61.430 -38.300 61.700 -38.030 ;
        RECT 68.180 -38.250 68.450 -37.980 ;
        RECT 74.930 -38.300 75.200 -38.030 ;
        RECT 81.680 -38.250 81.950 -37.980 ;
        RECT 88.430 -38.300 88.700 -38.030 ;
        RECT 95.180 -38.250 95.450 -37.980 ;
        RECT 101.930 -38.300 102.200 -38.030 ;
        RECT 108.680 -38.250 108.950 -37.980 ;
        RECT 115.430 -38.300 115.700 -38.030 ;
        RECT 122.180 -38.250 122.450 -37.980 ;
        RECT 128.930 -38.300 129.200 -38.030 ;
        RECT 135.680 -38.250 135.950 -37.980 ;
        RECT 142.430 -38.300 142.700 -38.030 ;
        RECT 149.180 -38.250 149.450 -37.980 ;
        RECT 155.930 -38.300 156.200 -38.030 ;
        RECT 162.680 -38.250 162.950 -37.980 ;
        RECT 169.430 -38.300 169.700 -38.030 ;
        RECT 176.180 -38.250 176.450 -37.980 ;
        RECT 182.930 -38.300 183.200 -38.030 ;
        RECT 189.680 -38.250 189.950 -37.980 ;
        RECT 196.430 -38.300 196.700 -38.030 ;
        RECT 203.180 -38.250 203.450 -37.980 ;
        RECT 209.930 -38.300 210.200 -38.030 ;
        RECT 216.680 -38.250 216.950 -37.980 ;
      LAYER met2 ;
        RECT 0.590 -37.890 1.070 -37.880 ;
        RECT 108.560 -37.890 109.070 -37.880 ;
        RECT 216.560 -37.890 217.040 -37.880 ;
        RECT 0.590 -38.410 217.040 -37.890 ;
    END
  END WL30
  PIN WL31
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER li1 ;
        RECT 0.590 -39.730 1.040 -39.290 ;
        RECT 14.090 -39.730 14.540 -39.290 ;
        RECT 27.590 -39.730 28.040 -39.290 ;
        RECT 41.090 -39.730 41.540 -39.290 ;
        RECT 54.590 -39.730 55.040 -39.290 ;
        RECT 68.090 -39.730 68.540 -39.290 ;
        RECT 81.590 -39.730 82.040 -39.290 ;
        RECT 95.090 -39.730 95.540 -39.290 ;
        RECT 108.590 -39.730 109.040 -39.290 ;
        RECT 122.090 -39.730 122.540 -39.290 ;
        RECT 135.590 -39.730 136.040 -39.290 ;
        RECT 149.090 -39.730 149.540 -39.290 ;
        RECT 162.590 -39.730 163.040 -39.290 ;
        RECT 176.090 -39.730 176.540 -39.290 ;
        RECT 189.590 -39.730 190.040 -39.290 ;
        RECT 203.090 -39.730 203.540 -39.290 ;
        RECT 216.590 -39.730 217.040 -39.290 ;
        RECT 7.340 -40.650 7.790 -40.200 ;
        RECT 20.840 -40.650 21.290 -40.200 ;
        RECT 34.340 -40.650 34.790 -40.200 ;
        RECT 47.840 -40.650 48.290 -40.200 ;
        RECT 61.340 -40.650 61.790 -40.200 ;
        RECT 74.840 -40.650 75.290 -40.200 ;
        RECT 88.340 -40.650 88.790 -40.200 ;
        RECT 101.840 -40.650 102.290 -40.200 ;
        RECT 115.340 -40.650 115.790 -40.200 ;
        RECT 128.840 -40.650 129.290 -40.200 ;
        RECT 142.340 -40.650 142.790 -40.200 ;
        RECT 155.840 -40.650 156.290 -40.200 ;
        RECT 169.340 -40.650 169.790 -40.200 ;
        RECT 182.840 -40.650 183.290 -40.200 ;
        RECT 196.340 -40.650 196.790 -40.200 ;
        RECT 209.840 -40.650 210.290 -40.200 ;
      LAYER mcon ;
        RECT 0.680 -39.650 0.950 -39.380 ;
        RECT 14.180 -39.650 14.450 -39.380 ;
        RECT 27.680 -39.650 27.950 -39.380 ;
        RECT 41.180 -39.650 41.450 -39.380 ;
        RECT 54.680 -39.650 54.950 -39.380 ;
        RECT 68.180 -39.650 68.450 -39.380 ;
        RECT 81.680 -39.650 81.950 -39.380 ;
        RECT 95.180 -39.650 95.450 -39.380 ;
        RECT 108.680 -39.650 108.950 -39.380 ;
        RECT 122.180 -39.650 122.450 -39.380 ;
        RECT 135.680 -39.650 135.950 -39.380 ;
        RECT 149.180 -39.650 149.450 -39.380 ;
        RECT 162.680 -39.650 162.950 -39.380 ;
        RECT 176.180 -39.650 176.450 -39.380 ;
        RECT 189.680 -39.650 189.950 -39.380 ;
        RECT 203.180 -39.650 203.450 -39.380 ;
        RECT 216.680 -39.650 216.950 -39.380 ;
        RECT 7.440 -40.550 7.690 -40.300 ;
        RECT 20.940 -40.550 21.190 -40.300 ;
        RECT 34.440 -40.550 34.690 -40.300 ;
        RECT 47.940 -40.550 48.190 -40.300 ;
        RECT 61.440 -40.550 61.690 -40.300 ;
        RECT 74.940 -40.550 75.190 -40.300 ;
        RECT 88.440 -40.550 88.690 -40.300 ;
        RECT 101.940 -40.550 102.190 -40.300 ;
        RECT 115.440 -40.550 115.690 -40.300 ;
        RECT 128.940 -40.550 129.190 -40.300 ;
        RECT 142.440 -40.550 142.690 -40.300 ;
        RECT 155.940 -40.550 156.190 -40.300 ;
        RECT 169.440 -40.550 169.690 -40.300 ;
        RECT 182.940 -40.550 183.190 -40.300 ;
        RECT 196.440 -40.550 196.690 -40.300 ;
        RECT 209.940 -40.550 210.190 -40.300 ;
      LAYER met1 ;
        RECT 0.580 -39.730 1.040 -39.290 ;
        RECT 0.580 -39.740 1.050 -39.730 ;
        RECT 0.590 -40.210 1.050 -39.740 ;
        RECT 7.330 -40.660 7.800 -39.730 ;
        RECT 14.080 -40.210 14.550 -39.290 ;
        RECT 20.830 -40.660 21.300 -39.730 ;
        RECT 27.580 -40.210 28.050 -39.290 ;
        RECT 34.330 -40.660 34.800 -39.730 ;
        RECT 41.080 -40.210 41.550 -39.290 ;
        RECT 47.830 -40.660 48.300 -39.730 ;
        RECT 54.580 -40.210 55.050 -39.290 ;
        RECT 61.330 -40.660 61.800 -39.730 ;
        RECT 68.080 -40.210 68.550 -39.290 ;
        RECT 74.830 -40.660 75.300 -39.730 ;
        RECT 81.580 -40.210 82.050 -39.290 ;
        RECT 88.330 -40.660 88.800 -39.730 ;
        RECT 95.080 -40.210 95.550 -39.290 ;
        RECT 101.830 -40.660 102.300 -39.730 ;
        RECT 108.580 -40.210 109.050 -39.290 ;
        RECT 115.330 -40.660 115.800 -39.730 ;
        RECT 122.080 -40.210 122.550 -39.290 ;
        RECT 128.830 -40.660 129.300 -39.730 ;
        RECT 135.580 -40.210 136.050 -39.290 ;
        RECT 142.330 -40.660 142.800 -39.730 ;
        RECT 149.080 -40.210 149.550 -39.290 ;
        RECT 155.830 -40.660 156.300 -39.730 ;
        RECT 162.580 -40.210 163.050 -39.290 ;
        RECT 169.330 -40.660 169.800 -39.730 ;
        RECT 176.080 -40.210 176.550 -39.290 ;
        RECT 182.830 -40.660 183.300 -39.730 ;
        RECT 189.580 -40.210 190.050 -39.290 ;
        RECT 196.330 -40.660 196.800 -39.730 ;
        RECT 203.080 -40.210 203.550 -39.290 ;
        RECT 216.590 -39.730 217.050 -39.290 ;
        RECT 209.830 -40.660 210.300 -39.730 ;
        RECT 216.580 -39.740 217.050 -39.730 ;
        RECT 216.580 -40.210 217.040 -39.740 ;
      LAYER via ;
        RECT 0.680 -40.150 0.950 -39.880 ;
        RECT 7.430 -40.130 7.700 -39.860 ;
        RECT 14.180 -40.150 14.450 -39.880 ;
        RECT 20.930 -40.130 21.200 -39.860 ;
        RECT 27.680 -40.150 27.950 -39.880 ;
        RECT 34.430 -40.130 34.700 -39.860 ;
        RECT 41.180 -40.150 41.450 -39.880 ;
        RECT 47.930 -40.130 48.200 -39.860 ;
        RECT 54.680 -40.150 54.950 -39.880 ;
        RECT 61.430 -40.130 61.700 -39.860 ;
        RECT 68.180 -40.150 68.450 -39.880 ;
        RECT 74.930 -40.130 75.200 -39.860 ;
        RECT 81.680 -40.150 81.950 -39.880 ;
        RECT 88.430 -40.130 88.700 -39.860 ;
        RECT 95.180 -40.150 95.450 -39.880 ;
        RECT 101.930 -40.130 102.200 -39.860 ;
        RECT 108.680 -40.150 108.950 -39.880 ;
        RECT 115.430 -40.130 115.700 -39.860 ;
        RECT 122.180 -40.150 122.450 -39.880 ;
        RECT 128.930 -40.130 129.200 -39.860 ;
        RECT 135.680 -40.150 135.950 -39.880 ;
        RECT 142.430 -40.130 142.700 -39.860 ;
        RECT 149.180 -40.150 149.450 -39.880 ;
        RECT 155.930 -40.130 156.200 -39.860 ;
        RECT 162.680 -40.150 162.950 -39.880 ;
        RECT 169.430 -40.130 169.700 -39.860 ;
        RECT 176.180 -40.150 176.450 -39.880 ;
        RECT 182.930 -40.130 183.200 -39.860 ;
        RECT 189.680 -40.150 189.950 -39.880 ;
        RECT 196.430 -40.130 196.700 -39.860 ;
        RECT 203.180 -40.150 203.450 -39.880 ;
        RECT 209.930 -40.130 210.200 -39.860 ;
        RECT 216.680 -40.150 216.950 -39.880 ;
      LAYER met2 ;
        RECT 0.590 -39.740 217.040 -39.730 ;
        RECT 0.580 -40.250 217.050 -39.740 ;
    END
  END WL31
  PIN BL16
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER li1 ;
        RECT 109.420 14.860 109.870 15.310 ;
        RECT 109.420 11.250 109.870 11.700 ;
        RECT 109.420 7.640 109.870 8.090 ;
        RECT 109.420 4.030 109.870 4.480 ;
        RECT 109.420 0.420 109.870 0.870 ;
        RECT 109.420 -3.190 109.870 -2.740 ;
        RECT 109.420 -6.800 109.870 -6.350 ;
        RECT 109.420 -10.410 109.870 -9.960 ;
        RECT 109.420 -14.020 109.870 -13.570 ;
        RECT 109.420 -17.630 109.870 -17.180 ;
        RECT 109.420 -21.240 109.870 -20.790 ;
        RECT 109.420 -24.850 109.870 -24.400 ;
        RECT 109.420 -28.460 109.870 -28.010 ;
        RECT 109.420 -32.070 109.870 -31.620 ;
        RECT 109.420 -35.680 109.870 -35.230 ;
        RECT 109.420 -39.290 109.870 -38.840 ;
      LAYER mcon ;
        RECT 109.520 14.960 109.770 15.210 ;
        RECT 109.520 11.350 109.770 11.600 ;
        RECT 109.520 7.740 109.770 7.990 ;
        RECT 109.520 4.130 109.770 4.380 ;
        RECT 109.520 0.520 109.770 0.770 ;
        RECT 109.520 -3.090 109.770 -2.840 ;
        RECT 109.520 -6.700 109.770 -6.450 ;
        RECT 109.520 -10.310 109.770 -10.060 ;
        RECT 109.520 -13.920 109.770 -13.670 ;
        RECT 109.520 -17.530 109.770 -17.280 ;
        RECT 109.520 -21.140 109.770 -20.890 ;
        RECT 109.520 -24.750 109.770 -24.500 ;
        RECT 109.520 -28.360 109.770 -28.110 ;
        RECT 109.520 -31.970 109.770 -31.720 ;
        RECT 109.520 -35.580 109.770 -35.330 ;
        RECT 109.520 -39.190 109.770 -38.940 ;
      LAYER met1 ;
        RECT 109.300 -43.100 109.980 19.120 ;
    END
  END BL16
  PIN BLb16
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER li1 ;
        RECT 114.520 16.660 114.970 17.110 ;
        RECT 114.520 13.050 114.970 13.510 ;
        RECT 114.520 9.440 114.970 9.900 ;
        RECT 114.520 5.830 114.970 6.290 ;
        RECT 114.520 2.220 114.970 2.680 ;
        RECT 114.520 -1.390 114.970 -0.930 ;
        RECT 114.520 -5.000 114.970 -4.540 ;
        RECT 114.520 -8.610 114.970 -8.150 ;
        RECT 114.520 -12.220 114.970 -11.760 ;
        RECT 114.520 -15.830 114.970 -15.370 ;
        RECT 114.520 -19.440 114.970 -18.980 ;
        RECT 114.520 -23.050 114.970 -22.590 ;
        RECT 114.520 -26.660 114.970 -26.200 ;
        RECT 114.520 -30.270 114.970 -29.810 ;
        RECT 114.520 -33.880 114.970 -33.420 ;
        RECT 114.520 -37.490 114.970 -37.030 ;
        RECT 114.520 -41.090 114.970 -40.640 ;
      LAYER mcon ;
        RECT 114.620 16.760 114.880 17.020 ;
        RECT 114.620 13.150 114.880 13.410 ;
        RECT 114.620 9.540 114.880 9.800 ;
        RECT 114.620 5.930 114.880 6.190 ;
        RECT 114.620 2.320 114.880 2.580 ;
        RECT 114.620 -1.290 114.880 -1.030 ;
        RECT 114.620 -4.900 114.880 -4.640 ;
        RECT 114.620 -8.510 114.880 -8.250 ;
        RECT 114.620 -12.120 114.880 -11.860 ;
        RECT 114.620 -15.730 114.880 -15.470 ;
        RECT 114.620 -19.340 114.880 -19.080 ;
        RECT 114.620 -22.950 114.880 -22.690 ;
        RECT 114.620 -26.560 114.880 -26.300 ;
        RECT 114.620 -30.170 114.880 -29.910 ;
        RECT 114.620 -33.780 114.880 -33.520 ;
        RECT 114.620 -37.390 114.880 -37.130 ;
        RECT 114.620 -41.000 114.880 -40.740 ;
      LAYER met1 ;
        RECT 114.400 -43.120 115.080 19.140 ;
    END
  END BLb16
  PIN BL17
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER li1 ;
        RECT 116.160 16.660 116.610 17.110 ;
        RECT 116.160 13.050 116.610 13.510 ;
        RECT 116.160 9.440 116.610 9.900 ;
        RECT 116.160 5.830 116.610 6.290 ;
        RECT 116.160 2.220 116.610 2.680 ;
        RECT 116.160 -1.390 116.610 -0.930 ;
        RECT 116.160 -5.000 116.610 -4.540 ;
        RECT 116.160 -8.610 116.610 -8.150 ;
        RECT 116.160 -12.220 116.610 -11.760 ;
        RECT 116.160 -15.830 116.610 -15.370 ;
        RECT 116.160 -19.440 116.610 -18.980 ;
        RECT 116.160 -23.050 116.610 -22.590 ;
        RECT 116.160 -26.660 116.610 -26.200 ;
        RECT 116.160 -30.270 116.610 -29.810 ;
        RECT 116.160 -33.880 116.610 -33.420 ;
        RECT 116.160 -37.490 116.610 -37.030 ;
        RECT 116.160 -41.090 116.610 -40.640 ;
      LAYER mcon ;
        RECT 116.250 16.760 116.510 17.020 ;
        RECT 116.250 13.150 116.510 13.410 ;
        RECT 116.250 9.540 116.510 9.800 ;
        RECT 116.250 5.930 116.510 6.190 ;
        RECT 116.250 2.320 116.510 2.580 ;
        RECT 116.250 -1.290 116.510 -1.030 ;
        RECT 116.250 -4.900 116.510 -4.640 ;
        RECT 116.250 -8.510 116.510 -8.250 ;
        RECT 116.250 -12.120 116.510 -11.860 ;
        RECT 116.250 -15.730 116.510 -15.470 ;
        RECT 116.250 -19.340 116.510 -19.080 ;
        RECT 116.250 -22.950 116.510 -22.690 ;
        RECT 116.250 -26.560 116.510 -26.300 ;
        RECT 116.250 -30.170 116.510 -29.910 ;
        RECT 116.250 -33.780 116.510 -33.520 ;
        RECT 116.250 -37.390 116.510 -37.130 ;
        RECT 116.250 -41.000 116.510 -40.740 ;
      LAYER met1 ;
        RECT 116.040 -43.110 116.720 19.130 ;
    END
  END BL17
  PIN BLb17
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER li1 ;
        RECT 121.260 14.860 121.710 15.310 ;
        RECT 121.260 11.250 121.710 11.700 ;
        RECT 121.260 7.640 121.710 8.090 ;
        RECT 121.260 4.030 121.710 4.480 ;
        RECT 121.260 0.420 121.710 0.870 ;
        RECT 121.260 -3.190 121.710 -2.740 ;
        RECT 121.260 -6.800 121.710 -6.350 ;
        RECT 121.260 -10.410 121.710 -9.960 ;
        RECT 121.260 -14.020 121.710 -13.570 ;
        RECT 121.260 -17.630 121.710 -17.180 ;
        RECT 121.260 -21.240 121.710 -20.790 ;
        RECT 121.260 -24.850 121.710 -24.400 ;
        RECT 121.260 -28.460 121.710 -28.010 ;
        RECT 121.260 -32.070 121.710 -31.620 ;
        RECT 121.260 -35.680 121.710 -35.230 ;
        RECT 121.260 -39.290 121.710 -38.840 ;
      LAYER mcon ;
        RECT 121.360 14.960 121.610 15.210 ;
        RECT 121.360 11.350 121.610 11.600 ;
        RECT 121.360 7.740 121.610 7.990 ;
        RECT 121.360 4.130 121.610 4.380 ;
        RECT 121.360 0.520 121.610 0.770 ;
        RECT 121.360 -3.090 121.610 -2.840 ;
        RECT 121.360 -6.700 121.610 -6.450 ;
        RECT 121.360 -10.310 121.610 -10.060 ;
        RECT 121.360 -13.920 121.610 -13.670 ;
        RECT 121.360 -17.530 121.610 -17.280 ;
        RECT 121.360 -21.140 121.610 -20.890 ;
        RECT 121.360 -24.750 121.610 -24.500 ;
        RECT 121.360 -28.360 121.610 -28.110 ;
        RECT 121.360 -31.970 121.610 -31.720 ;
        RECT 121.360 -35.580 121.610 -35.330 ;
        RECT 121.360 -39.190 121.610 -38.940 ;
      LAYER met1 ;
        RECT 121.160 -43.110 121.840 19.130 ;
    END
  END BLb17
  PIN BL18
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER li1 ;
        RECT 122.920 14.860 123.370 15.310 ;
        RECT 122.920 11.250 123.370 11.700 ;
        RECT 122.920 7.640 123.370 8.090 ;
        RECT 122.920 4.030 123.370 4.480 ;
        RECT 122.920 0.420 123.370 0.870 ;
        RECT 122.920 -3.190 123.370 -2.740 ;
        RECT 122.920 -6.800 123.370 -6.350 ;
        RECT 122.920 -10.410 123.370 -9.960 ;
        RECT 122.920 -14.020 123.370 -13.570 ;
        RECT 122.920 -17.630 123.370 -17.180 ;
        RECT 122.920 -21.240 123.370 -20.790 ;
        RECT 122.920 -24.850 123.370 -24.400 ;
        RECT 122.920 -28.460 123.370 -28.010 ;
        RECT 122.920 -32.070 123.370 -31.620 ;
        RECT 122.920 -35.680 123.370 -35.230 ;
        RECT 122.920 -39.290 123.370 -38.840 ;
      LAYER mcon ;
        RECT 123.020 14.960 123.270 15.210 ;
        RECT 123.020 11.350 123.270 11.600 ;
        RECT 123.020 7.740 123.270 7.990 ;
        RECT 123.020 4.130 123.270 4.380 ;
        RECT 123.020 0.520 123.270 0.770 ;
        RECT 123.020 -3.090 123.270 -2.840 ;
        RECT 123.020 -6.700 123.270 -6.450 ;
        RECT 123.020 -10.310 123.270 -10.060 ;
        RECT 123.020 -13.920 123.270 -13.670 ;
        RECT 123.020 -17.530 123.270 -17.280 ;
        RECT 123.020 -21.140 123.270 -20.890 ;
        RECT 123.020 -24.750 123.270 -24.500 ;
        RECT 123.020 -28.360 123.270 -28.110 ;
        RECT 123.020 -31.970 123.270 -31.720 ;
        RECT 123.020 -35.580 123.270 -35.330 ;
        RECT 123.020 -39.190 123.270 -38.940 ;
      LAYER met1 ;
        RECT 122.800 -43.110 123.480 19.130 ;
    END
  END BL18
  PIN BLb18
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER li1 ;
        RECT 128.020 16.660 128.470 17.110 ;
        RECT 128.020 13.050 128.470 13.510 ;
        RECT 128.020 9.440 128.470 9.900 ;
        RECT 128.020 5.830 128.470 6.290 ;
        RECT 128.020 2.220 128.470 2.680 ;
        RECT 128.020 -1.390 128.470 -0.930 ;
        RECT 128.020 -5.000 128.470 -4.540 ;
        RECT 128.020 -8.610 128.470 -8.150 ;
        RECT 128.020 -12.220 128.470 -11.760 ;
        RECT 128.020 -15.830 128.470 -15.370 ;
        RECT 128.020 -19.440 128.470 -18.980 ;
        RECT 128.020 -23.050 128.470 -22.590 ;
        RECT 128.020 -26.660 128.470 -26.200 ;
        RECT 128.020 -30.270 128.470 -29.810 ;
        RECT 128.020 -33.880 128.470 -33.420 ;
        RECT 128.020 -37.490 128.470 -37.030 ;
        RECT 128.020 -41.090 128.470 -40.640 ;
      LAYER mcon ;
        RECT 128.120 16.760 128.380 17.020 ;
        RECT 128.120 13.150 128.380 13.410 ;
        RECT 128.120 9.540 128.380 9.800 ;
        RECT 128.120 5.930 128.380 6.190 ;
        RECT 128.120 2.320 128.380 2.580 ;
        RECT 128.120 -1.290 128.380 -1.030 ;
        RECT 128.120 -4.900 128.380 -4.640 ;
        RECT 128.120 -8.510 128.380 -8.250 ;
        RECT 128.120 -12.120 128.380 -11.860 ;
        RECT 128.120 -15.730 128.380 -15.470 ;
        RECT 128.120 -19.340 128.380 -19.080 ;
        RECT 128.120 -22.950 128.380 -22.690 ;
        RECT 128.120 -26.560 128.380 -26.300 ;
        RECT 128.120 -30.170 128.380 -29.910 ;
        RECT 128.120 -33.780 128.380 -33.520 ;
        RECT 128.120 -37.390 128.380 -37.130 ;
        RECT 128.120 -41.000 128.380 -40.740 ;
      LAYER met1 ;
        RECT 127.910 -43.120 128.590 19.140 ;
    END
  END BLb18
  PIN BL19
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER li1 ;
        RECT 129.660 16.660 130.110 17.110 ;
        RECT 129.660 13.050 130.110 13.510 ;
        RECT 129.660 9.440 130.110 9.900 ;
        RECT 129.660 5.830 130.110 6.290 ;
        RECT 129.660 2.220 130.110 2.680 ;
        RECT 129.660 -1.390 130.110 -0.930 ;
        RECT 129.660 -5.000 130.110 -4.540 ;
        RECT 129.660 -8.610 130.110 -8.150 ;
        RECT 129.660 -12.220 130.110 -11.760 ;
        RECT 129.660 -15.830 130.110 -15.370 ;
        RECT 129.660 -19.440 130.110 -18.980 ;
        RECT 129.660 -23.050 130.110 -22.590 ;
        RECT 129.660 -26.660 130.110 -26.200 ;
        RECT 129.660 -30.270 130.110 -29.810 ;
        RECT 129.660 -33.880 130.110 -33.420 ;
        RECT 129.660 -37.490 130.110 -37.030 ;
        RECT 129.660 -41.090 130.110 -40.640 ;
      LAYER mcon ;
        RECT 129.750 16.760 130.010 17.020 ;
        RECT 129.750 13.150 130.010 13.410 ;
        RECT 129.750 9.540 130.010 9.800 ;
        RECT 129.750 5.930 130.010 6.190 ;
        RECT 129.750 2.320 130.010 2.580 ;
        RECT 129.750 -1.290 130.010 -1.030 ;
        RECT 129.750 -4.900 130.010 -4.640 ;
        RECT 129.750 -8.510 130.010 -8.250 ;
        RECT 129.750 -12.120 130.010 -11.860 ;
        RECT 129.750 -15.730 130.010 -15.470 ;
        RECT 129.750 -19.340 130.010 -19.080 ;
        RECT 129.750 -22.950 130.010 -22.690 ;
        RECT 129.750 -26.560 130.010 -26.300 ;
        RECT 129.750 -30.170 130.010 -29.910 ;
        RECT 129.750 -33.780 130.010 -33.520 ;
        RECT 129.750 -37.390 130.010 -37.130 ;
        RECT 129.750 -41.000 130.010 -40.740 ;
      LAYER met1 ;
        RECT 129.550 -43.110 130.230 19.130 ;
    END
  END BL19
  PIN BLb19
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER li1 ;
        RECT 134.760 14.860 135.210 15.310 ;
        RECT 134.760 11.250 135.210 11.700 ;
        RECT 134.760 7.640 135.210 8.090 ;
        RECT 134.760 4.030 135.210 4.480 ;
        RECT 134.760 0.420 135.210 0.870 ;
        RECT 134.760 -3.190 135.210 -2.740 ;
        RECT 134.760 -6.800 135.210 -6.350 ;
        RECT 134.760 -10.410 135.210 -9.960 ;
        RECT 134.760 -14.020 135.210 -13.570 ;
        RECT 134.760 -17.630 135.210 -17.180 ;
        RECT 134.760 -21.240 135.210 -20.790 ;
        RECT 134.760 -24.850 135.210 -24.400 ;
        RECT 134.760 -28.460 135.210 -28.010 ;
        RECT 134.760 -32.070 135.210 -31.620 ;
        RECT 134.760 -35.680 135.210 -35.230 ;
        RECT 134.760 -39.290 135.210 -38.840 ;
      LAYER mcon ;
        RECT 134.860 14.960 135.110 15.210 ;
        RECT 134.860 11.350 135.110 11.600 ;
        RECT 134.860 7.740 135.110 7.990 ;
        RECT 134.860 4.130 135.110 4.380 ;
        RECT 134.860 0.520 135.110 0.770 ;
        RECT 134.860 -3.090 135.110 -2.840 ;
        RECT 134.860 -6.700 135.110 -6.450 ;
        RECT 134.860 -10.310 135.110 -10.060 ;
        RECT 134.860 -13.920 135.110 -13.670 ;
        RECT 134.860 -17.530 135.110 -17.280 ;
        RECT 134.860 -21.140 135.110 -20.890 ;
        RECT 134.860 -24.750 135.110 -24.500 ;
        RECT 134.860 -28.360 135.110 -28.110 ;
        RECT 134.860 -31.970 135.110 -31.720 ;
        RECT 134.860 -35.580 135.110 -35.330 ;
        RECT 134.860 -39.190 135.110 -38.940 ;
      LAYER met1 ;
        RECT 134.650 -43.100 135.330 19.120 ;
    END
  END BLb19
  PIN BL20
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER li1 ;
        RECT 136.420 14.860 136.870 15.310 ;
        RECT 136.420 11.250 136.870 11.700 ;
        RECT 136.420 7.640 136.870 8.090 ;
        RECT 136.420 4.030 136.870 4.480 ;
        RECT 136.420 0.420 136.870 0.870 ;
        RECT 136.420 -3.190 136.870 -2.740 ;
        RECT 136.420 -6.800 136.870 -6.350 ;
        RECT 136.420 -10.410 136.870 -9.960 ;
        RECT 136.420 -14.020 136.870 -13.570 ;
        RECT 136.420 -17.630 136.870 -17.180 ;
        RECT 136.420 -21.240 136.870 -20.790 ;
        RECT 136.420 -24.850 136.870 -24.400 ;
        RECT 136.420 -28.460 136.870 -28.010 ;
        RECT 136.420 -32.070 136.870 -31.620 ;
        RECT 136.420 -35.680 136.870 -35.230 ;
        RECT 136.420 -39.290 136.870 -38.840 ;
      LAYER mcon ;
        RECT 136.520 14.960 136.770 15.210 ;
        RECT 136.520 11.350 136.770 11.600 ;
        RECT 136.520 7.740 136.770 7.990 ;
        RECT 136.520 4.130 136.770 4.380 ;
        RECT 136.520 0.520 136.770 0.770 ;
        RECT 136.520 -3.090 136.770 -2.840 ;
        RECT 136.520 -6.700 136.770 -6.450 ;
        RECT 136.520 -10.310 136.770 -10.060 ;
        RECT 136.520 -13.920 136.770 -13.670 ;
        RECT 136.520 -17.530 136.770 -17.280 ;
        RECT 136.520 -21.140 136.770 -20.890 ;
        RECT 136.520 -24.750 136.770 -24.500 ;
        RECT 136.520 -28.360 136.770 -28.110 ;
        RECT 136.520 -31.970 136.770 -31.720 ;
        RECT 136.520 -35.580 136.770 -35.330 ;
        RECT 136.520 -39.190 136.770 -38.940 ;
      LAYER met1 ;
        RECT 136.300 -43.100 136.980 19.120 ;
    END
  END BL20
  PIN BLb20
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER li1 ;
        RECT 141.520 16.660 141.970 17.110 ;
        RECT 141.520 13.050 141.970 13.510 ;
        RECT 141.520 9.440 141.970 9.900 ;
        RECT 141.520 5.830 141.970 6.290 ;
        RECT 141.520 2.220 141.970 2.680 ;
        RECT 141.520 -1.390 141.970 -0.930 ;
        RECT 141.520 -5.000 141.970 -4.540 ;
        RECT 141.520 -8.610 141.970 -8.150 ;
        RECT 141.520 -12.220 141.970 -11.760 ;
        RECT 141.520 -15.830 141.970 -15.370 ;
        RECT 141.520 -19.440 141.970 -18.980 ;
        RECT 141.520 -23.050 141.970 -22.590 ;
        RECT 141.520 -26.660 141.970 -26.200 ;
        RECT 141.520 -30.270 141.970 -29.810 ;
        RECT 141.520 -33.880 141.970 -33.420 ;
        RECT 141.520 -37.490 141.970 -37.030 ;
        RECT 141.520 -41.090 141.970 -40.640 ;
      LAYER mcon ;
        RECT 141.620 16.760 141.880 17.020 ;
        RECT 141.620 13.150 141.880 13.410 ;
        RECT 141.620 9.540 141.880 9.800 ;
        RECT 141.620 5.930 141.880 6.190 ;
        RECT 141.620 2.320 141.880 2.580 ;
        RECT 141.620 -1.290 141.880 -1.030 ;
        RECT 141.620 -4.900 141.880 -4.640 ;
        RECT 141.620 -8.510 141.880 -8.250 ;
        RECT 141.620 -12.120 141.880 -11.860 ;
        RECT 141.620 -15.730 141.880 -15.470 ;
        RECT 141.620 -19.340 141.880 -19.080 ;
        RECT 141.620 -22.950 141.880 -22.690 ;
        RECT 141.620 -26.560 141.880 -26.300 ;
        RECT 141.620 -30.170 141.880 -29.910 ;
        RECT 141.620 -33.780 141.880 -33.520 ;
        RECT 141.620 -37.390 141.880 -37.130 ;
        RECT 141.620 -41.000 141.880 -40.740 ;
      LAYER met1 ;
        RECT 141.400 -43.110 142.080 19.130 ;
    END
  END BLb20
  PIN BL21
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER li1 ;
        RECT 143.160 16.660 143.610 17.110 ;
        RECT 143.160 13.050 143.610 13.510 ;
        RECT 143.160 9.440 143.610 9.900 ;
        RECT 143.160 5.830 143.610 6.290 ;
        RECT 143.160 2.220 143.610 2.680 ;
        RECT 143.160 -1.390 143.610 -0.930 ;
        RECT 143.160 -5.000 143.610 -4.540 ;
        RECT 143.160 -8.610 143.610 -8.150 ;
        RECT 143.160 -12.220 143.610 -11.760 ;
        RECT 143.160 -15.830 143.610 -15.370 ;
        RECT 143.160 -19.440 143.610 -18.980 ;
        RECT 143.160 -23.050 143.610 -22.590 ;
        RECT 143.160 -26.660 143.610 -26.200 ;
        RECT 143.160 -30.270 143.610 -29.810 ;
        RECT 143.160 -33.880 143.610 -33.420 ;
        RECT 143.160 -37.490 143.610 -37.030 ;
        RECT 143.160 -41.090 143.610 -40.640 ;
      LAYER mcon ;
        RECT 143.250 16.760 143.510 17.020 ;
        RECT 143.250 13.150 143.510 13.410 ;
        RECT 143.250 9.540 143.510 9.800 ;
        RECT 143.250 5.930 143.510 6.190 ;
        RECT 143.250 2.320 143.510 2.580 ;
        RECT 143.250 -1.290 143.510 -1.030 ;
        RECT 143.250 -4.900 143.510 -4.640 ;
        RECT 143.250 -8.510 143.510 -8.250 ;
        RECT 143.250 -12.120 143.510 -11.860 ;
        RECT 143.250 -15.730 143.510 -15.470 ;
        RECT 143.250 -19.340 143.510 -19.080 ;
        RECT 143.250 -22.950 143.510 -22.690 ;
        RECT 143.250 -26.560 143.510 -26.300 ;
        RECT 143.250 -30.170 143.510 -29.910 ;
        RECT 143.250 -33.780 143.510 -33.520 ;
        RECT 143.250 -37.390 143.510 -37.130 ;
        RECT 143.250 -41.000 143.510 -40.740 ;
      LAYER met1 ;
        RECT 143.040 -43.120 143.720 19.140 ;
    END
  END BL21
  PIN BLb21
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER li1 ;
        RECT 148.260 14.860 148.710 15.310 ;
        RECT 148.260 11.250 148.710 11.700 ;
        RECT 148.260 7.640 148.710 8.090 ;
        RECT 148.260 4.030 148.710 4.480 ;
        RECT 148.260 0.420 148.710 0.870 ;
        RECT 148.260 -3.190 148.710 -2.740 ;
        RECT 148.260 -6.800 148.710 -6.350 ;
        RECT 148.260 -10.410 148.710 -9.960 ;
        RECT 148.260 -14.020 148.710 -13.570 ;
        RECT 148.260 -17.630 148.710 -17.180 ;
        RECT 148.260 -21.240 148.710 -20.790 ;
        RECT 148.260 -24.850 148.710 -24.400 ;
        RECT 148.260 -28.460 148.710 -28.010 ;
        RECT 148.260 -32.070 148.710 -31.620 ;
        RECT 148.260 -35.680 148.710 -35.230 ;
        RECT 148.260 -39.290 148.710 -38.840 ;
      LAYER mcon ;
        RECT 148.360 14.960 148.610 15.210 ;
        RECT 148.360 11.350 148.610 11.600 ;
        RECT 148.360 7.740 148.610 7.990 ;
        RECT 148.360 4.130 148.610 4.380 ;
        RECT 148.360 0.520 148.610 0.770 ;
        RECT 148.360 -3.090 148.610 -2.840 ;
        RECT 148.360 -6.700 148.610 -6.450 ;
        RECT 148.360 -10.310 148.610 -10.060 ;
        RECT 148.360 -13.920 148.610 -13.670 ;
        RECT 148.360 -17.530 148.610 -17.280 ;
        RECT 148.360 -21.140 148.610 -20.890 ;
        RECT 148.360 -24.750 148.610 -24.500 ;
        RECT 148.360 -28.360 148.610 -28.110 ;
        RECT 148.360 -31.970 148.610 -31.720 ;
        RECT 148.360 -35.580 148.610 -35.330 ;
        RECT 148.360 -39.190 148.610 -38.940 ;
      LAYER met1 ;
        RECT 148.150 -43.110 148.830 19.130 ;
    END
  END BLb21
  PIN BL22
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER li1 ;
        RECT 149.920 14.860 150.370 15.310 ;
        RECT 149.920 11.250 150.370 11.700 ;
        RECT 149.920 7.640 150.370 8.090 ;
        RECT 149.920 4.030 150.370 4.480 ;
        RECT 149.920 0.420 150.370 0.870 ;
        RECT 149.920 -3.190 150.370 -2.740 ;
        RECT 149.920 -6.800 150.370 -6.350 ;
        RECT 149.920 -10.410 150.370 -9.960 ;
        RECT 149.920 -14.020 150.370 -13.570 ;
        RECT 149.920 -17.630 150.370 -17.180 ;
        RECT 149.920 -21.240 150.370 -20.790 ;
        RECT 149.920 -24.850 150.370 -24.400 ;
        RECT 149.920 -28.460 150.370 -28.010 ;
        RECT 149.920 -32.070 150.370 -31.620 ;
        RECT 149.920 -35.680 150.370 -35.230 ;
        RECT 149.920 -39.290 150.370 -38.840 ;
      LAYER mcon ;
        RECT 150.020 14.960 150.270 15.210 ;
        RECT 150.020 11.350 150.270 11.600 ;
        RECT 150.020 7.740 150.270 7.990 ;
        RECT 150.020 4.130 150.270 4.380 ;
        RECT 150.020 0.520 150.270 0.770 ;
        RECT 150.020 -3.090 150.270 -2.840 ;
        RECT 150.020 -6.700 150.270 -6.450 ;
        RECT 150.020 -10.310 150.270 -10.060 ;
        RECT 150.020 -13.920 150.270 -13.670 ;
        RECT 150.020 -17.530 150.270 -17.280 ;
        RECT 150.020 -21.140 150.270 -20.890 ;
        RECT 150.020 -24.750 150.270 -24.500 ;
        RECT 150.020 -28.360 150.270 -28.110 ;
        RECT 150.020 -31.970 150.270 -31.720 ;
        RECT 150.020 -35.580 150.270 -35.330 ;
        RECT 150.020 -39.190 150.270 -38.940 ;
      LAYER met1 ;
        RECT 149.790 -43.110 150.470 19.130 ;
    END
  END BL22
  PIN BLb22
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER li1 ;
        RECT 155.020 16.660 155.470 17.110 ;
        RECT 155.020 13.050 155.470 13.510 ;
        RECT 155.020 9.440 155.470 9.900 ;
        RECT 155.020 5.830 155.470 6.290 ;
        RECT 155.020 2.220 155.470 2.680 ;
        RECT 155.020 -1.390 155.470 -0.930 ;
        RECT 155.020 -5.000 155.470 -4.540 ;
        RECT 155.020 -8.610 155.470 -8.150 ;
        RECT 155.020 -12.220 155.470 -11.760 ;
        RECT 155.020 -15.830 155.470 -15.370 ;
        RECT 155.020 -19.440 155.470 -18.980 ;
        RECT 155.020 -23.050 155.470 -22.590 ;
        RECT 155.020 -26.660 155.470 -26.200 ;
        RECT 155.020 -30.270 155.470 -29.810 ;
        RECT 155.020 -33.880 155.470 -33.420 ;
        RECT 155.020 -37.490 155.470 -37.030 ;
        RECT 155.020 -41.090 155.470 -40.640 ;
      LAYER mcon ;
        RECT 155.120 16.760 155.380 17.020 ;
        RECT 155.120 13.150 155.380 13.410 ;
        RECT 155.120 9.540 155.380 9.800 ;
        RECT 155.120 5.930 155.380 6.190 ;
        RECT 155.120 2.320 155.380 2.580 ;
        RECT 155.120 -1.290 155.380 -1.030 ;
        RECT 155.120 -4.900 155.380 -4.640 ;
        RECT 155.120 -8.510 155.380 -8.250 ;
        RECT 155.120 -12.120 155.380 -11.860 ;
        RECT 155.120 -15.730 155.380 -15.470 ;
        RECT 155.120 -19.340 155.380 -19.080 ;
        RECT 155.120 -22.950 155.380 -22.690 ;
        RECT 155.120 -26.560 155.380 -26.300 ;
        RECT 155.120 -30.170 155.380 -29.910 ;
        RECT 155.120 -33.780 155.380 -33.520 ;
        RECT 155.120 -37.390 155.380 -37.130 ;
        RECT 155.120 -41.000 155.380 -40.740 ;
      LAYER met1 ;
        RECT 154.910 -43.110 155.590 19.130 ;
    END
  END BLb22
  PIN BL23
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER li1 ;
        RECT 156.660 16.660 157.110 17.110 ;
        RECT 156.660 13.050 157.110 13.510 ;
        RECT 156.660 9.440 157.110 9.900 ;
        RECT 156.660 5.830 157.110 6.290 ;
        RECT 156.660 2.220 157.110 2.680 ;
        RECT 156.660 -1.390 157.110 -0.930 ;
        RECT 156.660 -5.000 157.110 -4.540 ;
        RECT 156.660 -8.610 157.110 -8.150 ;
        RECT 156.660 -12.220 157.110 -11.760 ;
        RECT 156.660 -15.830 157.110 -15.370 ;
        RECT 156.660 -19.440 157.110 -18.980 ;
        RECT 156.660 -23.050 157.110 -22.590 ;
        RECT 156.660 -26.660 157.110 -26.200 ;
        RECT 156.660 -30.270 157.110 -29.810 ;
        RECT 156.660 -33.880 157.110 -33.420 ;
        RECT 156.660 -37.490 157.110 -37.030 ;
        RECT 156.660 -41.090 157.110 -40.640 ;
      LAYER mcon ;
        RECT 156.750 16.760 157.010 17.020 ;
        RECT 156.750 13.150 157.010 13.410 ;
        RECT 156.750 9.540 157.010 9.800 ;
        RECT 156.750 5.930 157.010 6.190 ;
        RECT 156.750 2.320 157.010 2.580 ;
        RECT 156.750 -1.290 157.010 -1.030 ;
        RECT 156.750 -4.900 157.010 -4.640 ;
        RECT 156.750 -8.510 157.010 -8.250 ;
        RECT 156.750 -12.120 157.010 -11.860 ;
        RECT 156.750 -15.730 157.010 -15.470 ;
        RECT 156.750 -19.340 157.010 -19.080 ;
        RECT 156.750 -22.950 157.010 -22.690 ;
        RECT 156.750 -26.560 157.010 -26.300 ;
        RECT 156.750 -30.170 157.010 -29.910 ;
        RECT 156.750 -33.780 157.010 -33.520 ;
        RECT 156.750 -37.390 157.010 -37.130 ;
        RECT 156.750 -41.000 157.010 -40.740 ;
      LAYER met1 ;
        RECT 156.550 -43.120 157.230 19.140 ;
    END
  END BL23
  PIN BLb23
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER li1 ;
        RECT 161.760 14.860 162.210 15.310 ;
        RECT 161.760 11.250 162.210 11.700 ;
        RECT 161.760 7.640 162.210 8.090 ;
        RECT 161.760 4.030 162.210 4.480 ;
        RECT 161.760 0.420 162.210 0.870 ;
        RECT 161.760 -3.190 162.210 -2.740 ;
        RECT 161.760 -6.800 162.210 -6.350 ;
        RECT 161.760 -10.410 162.210 -9.960 ;
        RECT 161.760 -14.020 162.210 -13.570 ;
        RECT 161.760 -17.630 162.210 -17.180 ;
        RECT 161.760 -21.240 162.210 -20.790 ;
        RECT 161.760 -24.850 162.210 -24.400 ;
        RECT 161.760 -28.460 162.210 -28.010 ;
        RECT 161.760 -32.070 162.210 -31.620 ;
        RECT 161.760 -35.680 162.210 -35.230 ;
        RECT 161.760 -39.290 162.210 -38.840 ;
      LAYER mcon ;
        RECT 161.860 14.960 162.110 15.210 ;
        RECT 161.860 11.350 162.110 11.600 ;
        RECT 161.860 7.740 162.110 7.990 ;
        RECT 161.860 4.130 162.110 4.380 ;
        RECT 161.860 0.520 162.110 0.770 ;
        RECT 161.860 -3.090 162.110 -2.840 ;
        RECT 161.860 -6.700 162.110 -6.450 ;
        RECT 161.860 -10.310 162.110 -10.060 ;
        RECT 161.860 -13.920 162.110 -13.670 ;
        RECT 161.860 -17.530 162.110 -17.280 ;
        RECT 161.860 -21.140 162.110 -20.890 ;
        RECT 161.860 -24.750 162.110 -24.500 ;
        RECT 161.860 -28.360 162.110 -28.110 ;
        RECT 161.860 -31.970 162.110 -31.720 ;
        RECT 161.860 -35.580 162.110 -35.330 ;
        RECT 161.860 -39.190 162.110 -38.940 ;
      LAYER met1 ;
        RECT 161.650 -43.100 162.330 19.120 ;
    END
  END BLb23
  PIN BL24
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER li1 ;
        RECT 163.420 14.860 163.870 15.310 ;
        RECT 163.420 11.250 163.870 11.700 ;
        RECT 163.420 7.640 163.870 8.090 ;
        RECT 163.420 4.030 163.870 4.480 ;
        RECT 163.420 0.420 163.870 0.870 ;
        RECT 163.420 -3.190 163.870 -2.740 ;
        RECT 163.420 -6.800 163.870 -6.350 ;
        RECT 163.420 -10.410 163.870 -9.960 ;
        RECT 163.420 -14.020 163.870 -13.570 ;
        RECT 163.420 -17.630 163.870 -17.180 ;
        RECT 163.420 -21.240 163.870 -20.790 ;
        RECT 163.420 -24.850 163.870 -24.400 ;
        RECT 163.420 -28.460 163.870 -28.010 ;
        RECT 163.420 -32.070 163.870 -31.620 ;
        RECT 163.420 -35.680 163.870 -35.230 ;
        RECT 163.420 -39.290 163.870 -38.840 ;
      LAYER mcon ;
        RECT 163.520 14.960 163.770 15.210 ;
        RECT 163.520 11.350 163.770 11.600 ;
        RECT 163.520 7.740 163.770 7.990 ;
        RECT 163.520 4.130 163.770 4.380 ;
        RECT 163.520 0.520 163.770 0.770 ;
        RECT 163.520 -3.090 163.770 -2.840 ;
        RECT 163.520 -6.700 163.770 -6.450 ;
        RECT 163.520 -10.310 163.770 -10.060 ;
        RECT 163.520 -13.920 163.770 -13.670 ;
        RECT 163.520 -17.530 163.770 -17.280 ;
        RECT 163.520 -21.140 163.770 -20.890 ;
        RECT 163.520 -24.750 163.770 -24.500 ;
        RECT 163.520 -28.360 163.770 -28.110 ;
        RECT 163.520 -31.970 163.770 -31.720 ;
        RECT 163.520 -35.580 163.770 -35.330 ;
        RECT 163.520 -39.190 163.770 -38.940 ;
      LAYER met1 ;
        RECT 163.300 -43.100 163.980 19.120 ;
    END
  END BL24
  PIN BLb24
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER li1 ;
        RECT 168.520 16.660 168.970 17.110 ;
        RECT 168.520 13.050 168.970 13.510 ;
        RECT 168.520 9.440 168.970 9.900 ;
        RECT 168.520 5.830 168.970 6.290 ;
        RECT 168.520 2.220 168.970 2.680 ;
        RECT 168.520 -1.390 168.970 -0.930 ;
        RECT 168.520 -5.000 168.970 -4.540 ;
        RECT 168.520 -8.610 168.970 -8.150 ;
        RECT 168.520 -12.220 168.970 -11.760 ;
        RECT 168.520 -15.830 168.970 -15.370 ;
        RECT 168.520 -19.440 168.970 -18.980 ;
        RECT 168.520 -23.050 168.970 -22.590 ;
        RECT 168.520 -26.660 168.970 -26.200 ;
        RECT 168.520 -30.270 168.970 -29.810 ;
        RECT 168.520 -33.880 168.970 -33.420 ;
        RECT 168.520 -37.490 168.970 -37.030 ;
        RECT 168.520 -41.090 168.970 -40.640 ;
      LAYER mcon ;
        RECT 168.620 16.760 168.880 17.020 ;
        RECT 168.620 13.150 168.880 13.410 ;
        RECT 168.620 9.540 168.880 9.800 ;
        RECT 168.620 5.930 168.880 6.190 ;
        RECT 168.620 2.320 168.880 2.580 ;
        RECT 168.620 -1.290 168.880 -1.030 ;
        RECT 168.620 -4.900 168.880 -4.640 ;
        RECT 168.620 -8.510 168.880 -8.250 ;
        RECT 168.620 -12.120 168.880 -11.860 ;
        RECT 168.620 -15.730 168.880 -15.470 ;
        RECT 168.620 -19.340 168.880 -19.080 ;
        RECT 168.620 -22.950 168.880 -22.690 ;
        RECT 168.620 -26.560 168.880 -26.300 ;
        RECT 168.620 -30.170 168.880 -29.910 ;
        RECT 168.620 -33.780 168.880 -33.520 ;
        RECT 168.620 -37.390 168.880 -37.130 ;
        RECT 168.620 -41.000 168.880 -40.740 ;
      LAYER met1 ;
        RECT 168.400 -43.120 169.080 19.140 ;
    END
  END BLb24
  PIN BL25
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER li1 ;
        RECT 170.160 16.660 170.610 17.110 ;
        RECT 170.160 13.050 170.610 13.510 ;
        RECT 170.160 9.440 170.610 9.900 ;
        RECT 170.160 5.830 170.610 6.290 ;
        RECT 170.160 2.220 170.610 2.680 ;
        RECT 170.160 -1.390 170.610 -0.930 ;
        RECT 170.160 -5.000 170.610 -4.540 ;
        RECT 170.160 -8.610 170.610 -8.150 ;
        RECT 170.160 -12.220 170.610 -11.760 ;
        RECT 170.160 -15.830 170.610 -15.370 ;
        RECT 170.160 -19.440 170.610 -18.980 ;
        RECT 170.160 -23.050 170.610 -22.590 ;
        RECT 170.160 -26.660 170.610 -26.200 ;
        RECT 170.160 -30.270 170.610 -29.810 ;
        RECT 170.160 -33.880 170.610 -33.420 ;
        RECT 170.160 -37.490 170.610 -37.030 ;
        RECT 170.160 -41.090 170.610 -40.640 ;
      LAYER mcon ;
        RECT 170.250 16.760 170.510 17.020 ;
        RECT 170.250 13.150 170.510 13.410 ;
        RECT 170.250 9.540 170.510 9.800 ;
        RECT 170.250 5.930 170.510 6.190 ;
        RECT 170.250 2.320 170.510 2.580 ;
        RECT 170.250 -1.290 170.510 -1.030 ;
        RECT 170.250 -4.900 170.510 -4.640 ;
        RECT 170.250 -8.510 170.510 -8.250 ;
        RECT 170.250 -12.120 170.510 -11.860 ;
        RECT 170.250 -15.730 170.510 -15.470 ;
        RECT 170.250 -19.340 170.510 -19.080 ;
        RECT 170.250 -22.950 170.510 -22.690 ;
        RECT 170.250 -26.560 170.510 -26.300 ;
        RECT 170.250 -30.170 170.510 -29.910 ;
        RECT 170.250 -33.780 170.510 -33.520 ;
        RECT 170.250 -37.390 170.510 -37.130 ;
        RECT 170.250 -41.000 170.510 -40.740 ;
      LAYER met1 ;
        RECT 170.040 -43.110 170.720 19.130 ;
    END
  END BL25
  PIN BLb25
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER li1 ;
        RECT 175.260 14.860 175.710 15.310 ;
        RECT 175.260 11.250 175.710 11.700 ;
        RECT 175.260 7.640 175.710 8.090 ;
        RECT 175.260 4.030 175.710 4.480 ;
        RECT 175.260 0.420 175.710 0.870 ;
        RECT 175.260 -3.190 175.710 -2.740 ;
        RECT 175.260 -6.800 175.710 -6.350 ;
        RECT 175.260 -10.410 175.710 -9.960 ;
        RECT 175.260 -14.020 175.710 -13.570 ;
        RECT 175.260 -17.630 175.710 -17.180 ;
        RECT 175.260 -21.240 175.710 -20.790 ;
        RECT 175.260 -24.850 175.710 -24.400 ;
        RECT 175.260 -28.460 175.710 -28.010 ;
        RECT 175.260 -32.070 175.710 -31.620 ;
        RECT 175.260 -35.680 175.710 -35.230 ;
        RECT 175.260 -39.290 175.710 -38.840 ;
      LAYER mcon ;
        RECT 175.360 14.960 175.610 15.210 ;
        RECT 175.360 11.350 175.610 11.600 ;
        RECT 175.360 7.740 175.610 7.990 ;
        RECT 175.360 4.130 175.610 4.380 ;
        RECT 175.360 0.520 175.610 0.770 ;
        RECT 175.360 -3.090 175.610 -2.840 ;
        RECT 175.360 -6.700 175.610 -6.450 ;
        RECT 175.360 -10.310 175.610 -10.060 ;
        RECT 175.360 -13.920 175.610 -13.670 ;
        RECT 175.360 -17.530 175.610 -17.280 ;
        RECT 175.360 -21.140 175.610 -20.890 ;
        RECT 175.360 -24.750 175.610 -24.500 ;
        RECT 175.360 -28.360 175.610 -28.110 ;
        RECT 175.360 -31.970 175.610 -31.720 ;
        RECT 175.360 -35.580 175.610 -35.330 ;
        RECT 175.360 -39.190 175.610 -38.940 ;
      LAYER met1 ;
        RECT 175.160 -43.110 175.840 19.130 ;
    END
  END BLb25
  PIN BL26
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER li1 ;
        RECT 176.920 14.860 177.370 15.310 ;
        RECT 176.920 11.250 177.370 11.700 ;
        RECT 176.920 7.640 177.370 8.090 ;
        RECT 176.920 4.030 177.370 4.480 ;
        RECT 176.920 0.420 177.370 0.870 ;
        RECT 176.920 -3.190 177.370 -2.740 ;
        RECT 176.920 -6.800 177.370 -6.350 ;
        RECT 176.920 -10.410 177.370 -9.960 ;
        RECT 176.920 -14.020 177.370 -13.570 ;
        RECT 176.920 -17.630 177.370 -17.180 ;
        RECT 176.920 -21.240 177.370 -20.790 ;
        RECT 176.920 -24.850 177.370 -24.400 ;
        RECT 176.920 -28.460 177.370 -28.010 ;
        RECT 176.920 -32.070 177.370 -31.620 ;
        RECT 176.920 -35.680 177.370 -35.230 ;
        RECT 176.920 -39.290 177.370 -38.840 ;
      LAYER mcon ;
        RECT 177.020 14.960 177.270 15.210 ;
        RECT 177.020 11.350 177.270 11.600 ;
        RECT 177.020 7.740 177.270 7.990 ;
        RECT 177.020 4.130 177.270 4.380 ;
        RECT 177.020 0.520 177.270 0.770 ;
        RECT 177.020 -3.090 177.270 -2.840 ;
        RECT 177.020 -6.700 177.270 -6.450 ;
        RECT 177.020 -10.310 177.270 -10.060 ;
        RECT 177.020 -13.920 177.270 -13.670 ;
        RECT 177.020 -17.530 177.270 -17.280 ;
        RECT 177.020 -21.140 177.270 -20.890 ;
        RECT 177.020 -24.750 177.270 -24.500 ;
        RECT 177.020 -28.360 177.270 -28.110 ;
        RECT 177.020 -31.970 177.270 -31.720 ;
        RECT 177.020 -35.580 177.270 -35.330 ;
        RECT 177.020 -39.190 177.270 -38.940 ;
      LAYER met1 ;
        RECT 176.800 -43.110 177.480 19.130 ;
    END
  END BL26
  PIN BLb26
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER li1 ;
        RECT 182.020 16.660 182.470 17.110 ;
        RECT 182.020 13.050 182.470 13.510 ;
        RECT 182.020 9.440 182.470 9.900 ;
        RECT 182.020 5.830 182.470 6.290 ;
        RECT 182.020 2.220 182.470 2.680 ;
        RECT 182.020 -1.390 182.470 -0.930 ;
        RECT 182.020 -5.000 182.470 -4.540 ;
        RECT 182.020 -8.610 182.470 -8.150 ;
        RECT 182.020 -12.220 182.470 -11.760 ;
        RECT 182.020 -15.830 182.470 -15.370 ;
        RECT 182.020 -19.440 182.470 -18.980 ;
        RECT 182.020 -23.050 182.470 -22.590 ;
        RECT 182.020 -26.660 182.470 -26.200 ;
        RECT 182.020 -30.270 182.470 -29.810 ;
        RECT 182.020 -33.880 182.470 -33.420 ;
        RECT 182.020 -37.490 182.470 -37.030 ;
        RECT 182.020 -41.090 182.470 -40.640 ;
      LAYER mcon ;
        RECT 182.120 16.760 182.380 17.020 ;
        RECT 182.120 13.150 182.380 13.410 ;
        RECT 182.120 9.540 182.380 9.800 ;
        RECT 182.120 5.930 182.380 6.190 ;
        RECT 182.120 2.320 182.380 2.580 ;
        RECT 182.120 -1.290 182.380 -1.030 ;
        RECT 182.120 -4.900 182.380 -4.640 ;
        RECT 182.120 -8.510 182.380 -8.250 ;
        RECT 182.120 -12.120 182.380 -11.860 ;
        RECT 182.120 -15.730 182.380 -15.470 ;
        RECT 182.120 -19.340 182.380 -19.080 ;
        RECT 182.120 -22.950 182.380 -22.690 ;
        RECT 182.120 -26.560 182.380 -26.300 ;
        RECT 182.120 -30.170 182.380 -29.910 ;
        RECT 182.120 -33.780 182.380 -33.520 ;
        RECT 182.120 -37.390 182.380 -37.130 ;
        RECT 182.120 -41.000 182.380 -40.740 ;
      LAYER met1 ;
        RECT 181.910 -43.120 182.590 19.140 ;
    END
  END BLb26
  PIN BL27
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER li1 ;
        RECT 183.660 16.660 184.110 17.110 ;
        RECT 183.660 13.050 184.110 13.510 ;
        RECT 183.660 9.440 184.110 9.900 ;
        RECT 183.660 5.830 184.110 6.290 ;
        RECT 183.660 2.220 184.110 2.680 ;
        RECT 183.660 -1.390 184.110 -0.930 ;
        RECT 183.660 -5.000 184.110 -4.540 ;
        RECT 183.660 -8.610 184.110 -8.150 ;
        RECT 183.660 -12.220 184.110 -11.760 ;
        RECT 183.660 -15.830 184.110 -15.370 ;
        RECT 183.660 -19.440 184.110 -18.980 ;
        RECT 183.660 -23.050 184.110 -22.590 ;
        RECT 183.660 -26.660 184.110 -26.200 ;
        RECT 183.660 -30.270 184.110 -29.810 ;
        RECT 183.660 -33.880 184.110 -33.420 ;
        RECT 183.660 -37.490 184.110 -37.030 ;
        RECT 183.660 -41.090 184.110 -40.640 ;
      LAYER mcon ;
        RECT 183.750 16.760 184.010 17.020 ;
        RECT 183.750 13.150 184.010 13.410 ;
        RECT 183.750 9.540 184.010 9.800 ;
        RECT 183.750 5.930 184.010 6.190 ;
        RECT 183.750 2.320 184.010 2.580 ;
        RECT 183.750 -1.290 184.010 -1.030 ;
        RECT 183.750 -4.900 184.010 -4.640 ;
        RECT 183.750 -8.510 184.010 -8.250 ;
        RECT 183.750 -12.120 184.010 -11.860 ;
        RECT 183.750 -15.730 184.010 -15.470 ;
        RECT 183.750 -19.340 184.010 -19.080 ;
        RECT 183.750 -22.950 184.010 -22.690 ;
        RECT 183.750 -26.560 184.010 -26.300 ;
        RECT 183.750 -30.170 184.010 -29.910 ;
        RECT 183.750 -33.780 184.010 -33.520 ;
        RECT 183.750 -37.390 184.010 -37.130 ;
        RECT 183.750 -41.000 184.010 -40.740 ;
      LAYER met1 ;
        RECT 183.550 -43.110 184.230 19.130 ;
    END
  END BL27
  PIN BLb27
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER li1 ;
        RECT 188.760 14.860 189.210 15.310 ;
        RECT 188.760 11.250 189.210 11.700 ;
        RECT 188.760 7.640 189.210 8.090 ;
        RECT 188.760 4.030 189.210 4.480 ;
        RECT 188.760 0.420 189.210 0.870 ;
        RECT 188.760 -3.190 189.210 -2.740 ;
        RECT 188.760 -6.800 189.210 -6.350 ;
        RECT 188.760 -10.410 189.210 -9.960 ;
        RECT 188.760 -14.020 189.210 -13.570 ;
        RECT 188.760 -17.630 189.210 -17.180 ;
        RECT 188.760 -21.240 189.210 -20.790 ;
        RECT 188.760 -24.850 189.210 -24.400 ;
        RECT 188.760 -28.460 189.210 -28.010 ;
        RECT 188.760 -32.070 189.210 -31.620 ;
        RECT 188.760 -35.680 189.210 -35.230 ;
        RECT 188.760 -39.290 189.210 -38.840 ;
      LAYER mcon ;
        RECT 188.860 14.960 189.110 15.210 ;
        RECT 188.860 11.350 189.110 11.600 ;
        RECT 188.860 7.740 189.110 7.990 ;
        RECT 188.860 4.130 189.110 4.380 ;
        RECT 188.860 0.520 189.110 0.770 ;
        RECT 188.860 -3.090 189.110 -2.840 ;
        RECT 188.860 -6.700 189.110 -6.450 ;
        RECT 188.860 -10.310 189.110 -10.060 ;
        RECT 188.860 -13.920 189.110 -13.670 ;
        RECT 188.860 -17.530 189.110 -17.280 ;
        RECT 188.860 -21.140 189.110 -20.890 ;
        RECT 188.860 -24.750 189.110 -24.500 ;
        RECT 188.860 -28.360 189.110 -28.110 ;
        RECT 188.860 -31.970 189.110 -31.720 ;
        RECT 188.860 -35.580 189.110 -35.330 ;
        RECT 188.860 -39.190 189.110 -38.940 ;
      LAYER met1 ;
        RECT 188.650 -43.100 189.330 19.120 ;
    END
  END BLb27
  PIN BL28
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER li1 ;
        RECT 190.420 14.860 190.870 15.310 ;
        RECT 190.420 11.250 190.870 11.700 ;
        RECT 190.420 7.640 190.870 8.090 ;
        RECT 190.420 4.030 190.870 4.480 ;
        RECT 190.420 0.420 190.870 0.870 ;
        RECT 190.420 -3.190 190.870 -2.740 ;
        RECT 190.420 -6.800 190.870 -6.350 ;
        RECT 190.420 -10.410 190.870 -9.960 ;
        RECT 190.420 -14.020 190.870 -13.570 ;
        RECT 190.420 -17.630 190.870 -17.180 ;
        RECT 190.420 -21.240 190.870 -20.790 ;
        RECT 190.420 -24.850 190.870 -24.400 ;
        RECT 190.420 -28.460 190.870 -28.010 ;
        RECT 190.420 -32.070 190.870 -31.620 ;
        RECT 190.420 -35.680 190.870 -35.230 ;
        RECT 190.420 -39.290 190.870 -38.840 ;
      LAYER mcon ;
        RECT 190.520 14.960 190.770 15.210 ;
        RECT 190.520 11.350 190.770 11.600 ;
        RECT 190.520 7.740 190.770 7.990 ;
        RECT 190.520 4.130 190.770 4.380 ;
        RECT 190.520 0.520 190.770 0.770 ;
        RECT 190.520 -3.090 190.770 -2.840 ;
        RECT 190.520 -6.700 190.770 -6.450 ;
        RECT 190.520 -10.310 190.770 -10.060 ;
        RECT 190.520 -13.920 190.770 -13.670 ;
        RECT 190.520 -17.530 190.770 -17.280 ;
        RECT 190.520 -21.140 190.770 -20.890 ;
        RECT 190.520 -24.750 190.770 -24.500 ;
        RECT 190.520 -28.360 190.770 -28.110 ;
        RECT 190.520 -31.970 190.770 -31.720 ;
        RECT 190.520 -35.580 190.770 -35.330 ;
        RECT 190.520 -39.190 190.770 -38.940 ;
      LAYER met1 ;
        RECT 190.300 -43.100 190.980 19.120 ;
    END
  END BL28
  PIN BLb28
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER li1 ;
        RECT 195.520 16.660 195.970 17.110 ;
        RECT 195.520 13.050 195.970 13.510 ;
        RECT 195.520 9.440 195.970 9.900 ;
        RECT 195.520 5.830 195.970 6.290 ;
        RECT 195.520 2.220 195.970 2.680 ;
        RECT 195.520 -1.390 195.970 -0.930 ;
        RECT 195.520 -5.000 195.970 -4.540 ;
        RECT 195.520 -8.610 195.970 -8.150 ;
        RECT 195.520 -12.220 195.970 -11.760 ;
        RECT 195.520 -15.830 195.970 -15.370 ;
        RECT 195.520 -19.440 195.970 -18.980 ;
        RECT 195.520 -23.050 195.970 -22.590 ;
        RECT 195.520 -26.660 195.970 -26.200 ;
        RECT 195.520 -30.270 195.970 -29.810 ;
        RECT 195.520 -33.880 195.970 -33.420 ;
        RECT 195.520 -37.490 195.970 -37.030 ;
        RECT 195.520 -41.090 195.970 -40.640 ;
      LAYER mcon ;
        RECT 195.620 16.760 195.880 17.020 ;
        RECT 195.620 13.150 195.880 13.410 ;
        RECT 195.620 9.540 195.880 9.800 ;
        RECT 195.620 5.930 195.880 6.190 ;
        RECT 195.620 2.320 195.880 2.580 ;
        RECT 195.620 -1.290 195.880 -1.030 ;
        RECT 195.620 -4.900 195.880 -4.640 ;
        RECT 195.620 -8.510 195.880 -8.250 ;
        RECT 195.620 -12.120 195.880 -11.860 ;
        RECT 195.620 -15.730 195.880 -15.470 ;
        RECT 195.620 -19.340 195.880 -19.080 ;
        RECT 195.620 -22.950 195.880 -22.690 ;
        RECT 195.620 -26.560 195.880 -26.300 ;
        RECT 195.620 -30.170 195.880 -29.910 ;
        RECT 195.620 -33.780 195.880 -33.520 ;
        RECT 195.620 -37.390 195.880 -37.130 ;
        RECT 195.620 -41.000 195.880 -40.740 ;
      LAYER met1 ;
        RECT 195.400 -43.110 196.080 19.130 ;
    END
  END BLb28
  PIN BL29
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER li1 ;
        RECT 197.160 16.660 197.610 17.110 ;
        RECT 197.160 13.050 197.610 13.510 ;
        RECT 197.160 9.440 197.610 9.900 ;
        RECT 197.160 5.830 197.610 6.290 ;
        RECT 197.160 2.220 197.610 2.680 ;
        RECT 197.160 -1.390 197.610 -0.930 ;
        RECT 197.160 -5.000 197.610 -4.540 ;
        RECT 197.160 -8.610 197.610 -8.150 ;
        RECT 197.160 -12.220 197.610 -11.760 ;
        RECT 197.160 -15.830 197.610 -15.370 ;
        RECT 197.160 -19.440 197.610 -18.980 ;
        RECT 197.160 -23.050 197.610 -22.590 ;
        RECT 197.160 -26.660 197.610 -26.200 ;
        RECT 197.160 -30.270 197.610 -29.810 ;
        RECT 197.160 -33.880 197.610 -33.420 ;
        RECT 197.160 -37.490 197.610 -37.030 ;
        RECT 197.160 -41.090 197.610 -40.640 ;
      LAYER mcon ;
        RECT 197.250 16.760 197.510 17.020 ;
        RECT 197.250 13.150 197.510 13.410 ;
        RECT 197.250 9.540 197.510 9.800 ;
        RECT 197.250 5.930 197.510 6.190 ;
        RECT 197.250 2.320 197.510 2.580 ;
        RECT 197.250 -1.290 197.510 -1.030 ;
        RECT 197.250 -4.900 197.510 -4.640 ;
        RECT 197.250 -8.510 197.510 -8.250 ;
        RECT 197.250 -12.120 197.510 -11.860 ;
        RECT 197.250 -15.730 197.510 -15.470 ;
        RECT 197.250 -19.340 197.510 -19.080 ;
        RECT 197.250 -22.950 197.510 -22.690 ;
        RECT 197.250 -26.560 197.510 -26.300 ;
        RECT 197.250 -30.170 197.510 -29.910 ;
        RECT 197.250 -33.780 197.510 -33.520 ;
        RECT 197.250 -37.390 197.510 -37.130 ;
        RECT 197.250 -41.000 197.510 -40.740 ;
      LAYER met1 ;
        RECT 197.040 -43.120 197.720 19.140 ;
    END
  END BL29
  PIN BLb29
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER li1 ;
        RECT 202.260 14.860 202.710 15.310 ;
        RECT 202.260 11.250 202.710 11.700 ;
        RECT 202.260 7.640 202.710 8.090 ;
        RECT 202.260 4.030 202.710 4.480 ;
        RECT 202.260 0.420 202.710 0.870 ;
        RECT 202.260 -3.190 202.710 -2.740 ;
        RECT 202.260 -6.800 202.710 -6.350 ;
        RECT 202.260 -10.410 202.710 -9.960 ;
        RECT 202.260 -14.020 202.710 -13.570 ;
        RECT 202.260 -17.630 202.710 -17.180 ;
        RECT 202.260 -21.240 202.710 -20.790 ;
        RECT 202.260 -24.850 202.710 -24.400 ;
        RECT 202.260 -28.460 202.710 -28.010 ;
        RECT 202.260 -32.070 202.710 -31.620 ;
        RECT 202.260 -35.680 202.710 -35.230 ;
        RECT 202.260 -39.290 202.710 -38.840 ;
      LAYER mcon ;
        RECT 202.360 14.960 202.610 15.210 ;
        RECT 202.360 11.350 202.610 11.600 ;
        RECT 202.360 7.740 202.610 7.990 ;
        RECT 202.360 4.130 202.610 4.380 ;
        RECT 202.360 0.520 202.610 0.770 ;
        RECT 202.360 -3.090 202.610 -2.840 ;
        RECT 202.360 -6.700 202.610 -6.450 ;
        RECT 202.360 -10.310 202.610 -10.060 ;
        RECT 202.360 -13.920 202.610 -13.670 ;
        RECT 202.360 -17.530 202.610 -17.280 ;
        RECT 202.360 -21.140 202.610 -20.890 ;
        RECT 202.360 -24.750 202.610 -24.500 ;
        RECT 202.360 -28.360 202.610 -28.110 ;
        RECT 202.360 -31.970 202.610 -31.720 ;
        RECT 202.360 -35.580 202.610 -35.330 ;
        RECT 202.360 -39.190 202.610 -38.940 ;
      LAYER met1 ;
        RECT 202.150 -43.110 202.830 19.130 ;
    END
  END BLb29
  PIN BL30
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER li1 ;
        RECT 203.920 14.860 204.370 15.310 ;
        RECT 203.920 11.250 204.370 11.700 ;
        RECT 203.920 7.640 204.370 8.090 ;
        RECT 203.920 4.030 204.370 4.480 ;
        RECT 203.920 0.420 204.370 0.870 ;
        RECT 203.920 -3.190 204.370 -2.740 ;
        RECT 203.920 -6.800 204.370 -6.350 ;
        RECT 203.920 -10.410 204.370 -9.960 ;
        RECT 203.920 -14.020 204.370 -13.570 ;
        RECT 203.920 -17.630 204.370 -17.180 ;
        RECT 203.920 -21.240 204.370 -20.790 ;
        RECT 203.920 -24.850 204.370 -24.400 ;
        RECT 203.920 -28.460 204.370 -28.010 ;
        RECT 203.920 -32.070 204.370 -31.620 ;
        RECT 203.920 -35.680 204.370 -35.230 ;
        RECT 203.920 -39.290 204.370 -38.840 ;
      LAYER mcon ;
        RECT 204.020 14.960 204.270 15.210 ;
        RECT 204.020 11.350 204.270 11.600 ;
        RECT 204.020 7.740 204.270 7.990 ;
        RECT 204.020 4.130 204.270 4.380 ;
        RECT 204.020 0.520 204.270 0.770 ;
        RECT 204.020 -3.090 204.270 -2.840 ;
        RECT 204.020 -6.700 204.270 -6.450 ;
        RECT 204.020 -10.310 204.270 -10.060 ;
        RECT 204.020 -13.920 204.270 -13.670 ;
        RECT 204.020 -17.530 204.270 -17.280 ;
        RECT 204.020 -21.140 204.270 -20.890 ;
        RECT 204.020 -24.750 204.270 -24.500 ;
        RECT 204.020 -28.360 204.270 -28.110 ;
        RECT 204.020 -31.970 204.270 -31.720 ;
        RECT 204.020 -35.580 204.270 -35.330 ;
        RECT 204.020 -39.190 204.270 -38.940 ;
      LAYER met1 ;
        RECT 203.790 -43.110 204.470 19.130 ;
    END
  END BL30
  PIN BLb30
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER li1 ;
        RECT 209.020 16.660 209.470 17.110 ;
        RECT 209.020 13.050 209.470 13.510 ;
        RECT 209.020 9.440 209.470 9.900 ;
        RECT 209.020 5.830 209.470 6.290 ;
        RECT 209.020 2.220 209.470 2.680 ;
        RECT 209.020 -1.390 209.470 -0.930 ;
        RECT 209.020 -5.000 209.470 -4.540 ;
        RECT 209.020 -8.610 209.470 -8.150 ;
        RECT 209.020 -12.220 209.470 -11.760 ;
        RECT 209.020 -15.830 209.470 -15.370 ;
        RECT 209.020 -19.440 209.470 -18.980 ;
        RECT 209.020 -23.050 209.470 -22.590 ;
        RECT 209.020 -26.660 209.470 -26.200 ;
        RECT 209.020 -30.270 209.470 -29.810 ;
        RECT 209.020 -33.880 209.470 -33.420 ;
        RECT 209.020 -37.490 209.470 -37.030 ;
        RECT 209.020 -41.090 209.470 -40.640 ;
      LAYER mcon ;
        RECT 209.120 16.760 209.380 17.020 ;
        RECT 209.120 13.150 209.380 13.410 ;
        RECT 209.120 9.540 209.380 9.800 ;
        RECT 209.120 5.930 209.380 6.190 ;
        RECT 209.120 2.320 209.380 2.580 ;
        RECT 209.120 -1.290 209.380 -1.030 ;
        RECT 209.120 -4.900 209.380 -4.640 ;
        RECT 209.120 -8.510 209.380 -8.250 ;
        RECT 209.120 -12.120 209.380 -11.860 ;
        RECT 209.120 -15.730 209.380 -15.470 ;
        RECT 209.120 -19.340 209.380 -19.080 ;
        RECT 209.120 -22.950 209.380 -22.690 ;
        RECT 209.120 -26.560 209.380 -26.300 ;
        RECT 209.120 -30.170 209.380 -29.910 ;
        RECT 209.120 -33.780 209.380 -33.520 ;
        RECT 209.120 -37.390 209.380 -37.130 ;
        RECT 209.120 -41.000 209.380 -40.740 ;
      LAYER met1 ;
        RECT 208.910 -43.110 209.590 19.130 ;
    END
  END BLb30
  PIN BL31
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER li1 ;
        RECT 210.660 16.660 211.110 17.110 ;
        RECT 210.660 13.050 211.110 13.510 ;
        RECT 210.660 9.440 211.110 9.900 ;
        RECT 210.660 5.830 211.110 6.290 ;
        RECT 210.660 2.220 211.110 2.680 ;
        RECT 210.660 -1.390 211.110 -0.930 ;
        RECT 210.660 -5.000 211.110 -4.540 ;
        RECT 210.660 -8.610 211.110 -8.150 ;
        RECT 210.660 -12.220 211.110 -11.760 ;
        RECT 210.660 -15.830 211.110 -15.370 ;
        RECT 210.660 -19.440 211.110 -18.980 ;
        RECT 210.660 -23.050 211.110 -22.590 ;
        RECT 210.660 -26.660 211.110 -26.200 ;
        RECT 210.660 -30.270 211.110 -29.810 ;
        RECT 210.660 -33.880 211.110 -33.420 ;
        RECT 210.660 -37.490 211.110 -37.030 ;
        RECT 210.660 -41.090 211.110 -40.640 ;
      LAYER mcon ;
        RECT 210.750 16.760 211.010 17.020 ;
        RECT 210.750 13.150 211.010 13.410 ;
        RECT 210.750 9.540 211.010 9.800 ;
        RECT 210.750 5.930 211.010 6.190 ;
        RECT 210.750 2.320 211.010 2.580 ;
        RECT 210.750 -1.290 211.010 -1.030 ;
        RECT 210.750 -4.900 211.010 -4.640 ;
        RECT 210.750 -8.510 211.010 -8.250 ;
        RECT 210.750 -12.120 211.010 -11.860 ;
        RECT 210.750 -15.730 211.010 -15.470 ;
        RECT 210.750 -19.340 211.010 -19.080 ;
        RECT 210.750 -22.950 211.010 -22.690 ;
        RECT 210.750 -26.560 211.010 -26.300 ;
        RECT 210.750 -30.170 211.010 -29.910 ;
        RECT 210.750 -33.780 211.010 -33.520 ;
        RECT 210.750 -37.390 211.010 -37.130 ;
        RECT 210.750 -41.000 211.010 -40.740 ;
      LAYER met1 ;
        RECT 210.550 -43.120 211.230 19.140 ;
    END
  END BL31
  PIN BLb31
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER li1 ;
        RECT 215.760 14.860 216.210 15.310 ;
        RECT 215.760 11.250 216.210 11.700 ;
        RECT 215.760 7.640 216.210 8.090 ;
        RECT 215.760 4.030 216.210 4.480 ;
        RECT 215.760 0.420 216.210 0.870 ;
        RECT 215.760 -3.190 216.210 -2.740 ;
        RECT 215.760 -6.800 216.210 -6.350 ;
        RECT 215.760 -10.410 216.210 -9.960 ;
        RECT 215.760 -14.020 216.210 -13.570 ;
        RECT 215.760 -17.630 216.210 -17.180 ;
        RECT 215.760 -21.240 216.210 -20.790 ;
        RECT 215.760 -24.850 216.210 -24.400 ;
        RECT 215.760 -28.460 216.210 -28.010 ;
        RECT 215.760 -32.070 216.210 -31.620 ;
        RECT 215.760 -35.680 216.210 -35.230 ;
        RECT 215.760 -39.290 216.210 -38.840 ;
      LAYER mcon ;
        RECT 215.860 14.960 216.110 15.210 ;
        RECT 215.860 11.350 216.110 11.600 ;
        RECT 215.860 7.740 216.110 7.990 ;
        RECT 215.860 4.130 216.110 4.380 ;
        RECT 215.860 0.520 216.110 0.770 ;
        RECT 215.860 -3.090 216.110 -2.840 ;
        RECT 215.860 -6.700 216.110 -6.450 ;
        RECT 215.860 -10.310 216.110 -10.060 ;
        RECT 215.860 -13.920 216.110 -13.670 ;
        RECT 215.860 -17.530 216.110 -17.280 ;
        RECT 215.860 -21.140 216.110 -20.890 ;
        RECT 215.860 -24.750 216.110 -24.500 ;
        RECT 215.860 -28.360 216.110 -28.110 ;
        RECT 215.860 -31.970 216.110 -31.720 ;
        RECT 215.860 -35.580 216.110 -35.330 ;
        RECT 215.860 -39.190 216.110 -38.940 ;
      LAYER met1 ;
        RECT 215.650 -43.100 216.330 19.120 ;
    END
  END BLb31
  PIN vccd1
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 2.970 -41.390 5.420 17.410 ;
        RECT 9.710 -41.390 12.160 17.410 ;
        RECT 16.470 -41.390 18.920 17.410 ;
        RECT 23.210 -41.390 25.660 17.410 ;
        RECT 29.970 -41.390 32.420 17.410 ;
        RECT 36.710 -41.390 39.160 17.410 ;
        RECT 43.470 -41.390 45.920 17.410 ;
        RECT 50.210 -41.390 52.660 17.410 ;
        RECT 56.970 -41.390 59.420 17.410 ;
        RECT 63.710 -41.390 66.160 17.410 ;
        RECT 70.470 -41.390 72.920 17.410 ;
        RECT 77.210 -41.390 79.660 17.410 ;
        RECT 83.970 -41.390 86.420 17.410 ;
        RECT 90.710 -41.390 93.160 17.410 ;
        RECT 97.470 -41.390 99.920 17.410 ;
        RECT 104.210 -41.390 106.660 17.410 ;
        RECT 110.970 -41.390 113.420 17.410 ;
        RECT 117.710 -41.390 120.160 17.410 ;
        RECT 124.470 -41.390 126.920 17.410 ;
        RECT 131.210 -41.390 133.660 17.410 ;
        RECT 137.970 -41.390 140.420 17.410 ;
        RECT 144.710 -41.390 147.160 17.410 ;
        RECT 151.470 -41.390 153.920 17.410 ;
        RECT 158.210 -41.390 160.660 17.410 ;
        RECT 164.970 -41.390 167.420 17.410 ;
        RECT 171.710 -41.390 174.160 17.410 ;
        RECT 178.470 -41.390 180.920 17.410 ;
        RECT 185.210 -41.390 187.660 17.410 ;
        RECT 191.970 -41.390 194.420 17.410 ;
        RECT 198.710 -41.390 201.160 17.410 ;
        RECT 205.470 -41.390 207.920 17.410 ;
        RECT 212.210 -41.390 214.660 17.410 ;
      LAYER li1 ;
        RECT 3.270 16.960 3.720 17.110 ;
        RECT 3.970 17.000 4.420 17.110 ;
        RECT 4.670 17.000 5.080 17.100 ;
        RECT 3.970 16.960 5.080 17.000 ;
        RECT 3.270 16.740 5.080 16.960 ;
        RECT 3.270 16.660 4.420 16.740 ;
        RECT 4.670 16.680 5.080 16.740 ;
        RECT 10.050 17.000 10.460 17.100 ;
        RECT 10.710 17.000 11.160 17.110 ;
        RECT 10.050 16.960 11.160 17.000 ;
        RECT 11.410 16.960 11.860 17.110 ;
        RECT 10.050 16.740 11.860 16.960 ;
        RECT 10.050 16.680 10.460 16.740 ;
        RECT 3.970 16.560 4.420 16.660 ;
        RECT 10.710 16.660 11.860 16.740 ;
        RECT 16.770 16.960 17.220 17.110 ;
        RECT 17.470 17.000 17.920 17.110 ;
        RECT 18.170 17.000 18.580 17.100 ;
        RECT 17.470 16.960 18.580 17.000 ;
        RECT 16.770 16.740 18.580 16.960 ;
        RECT 16.770 16.660 17.920 16.740 ;
        RECT 18.170 16.680 18.580 16.740 ;
        RECT 23.550 17.000 23.960 17.100 ;
        RECT 24.210 17.000 24.660 17.110 ;
        RECT 23.550 16.960 24.660 17.000 ;
        RECT 24.910 16.960 25.360 17.110 ;
        RECT 23.550 16.740 25.360 16.960 ;
        RECT 23.550 16.680 23.960 16.740 ;
        RECT 10.710 16.560 11.160 16.660 ;
        RECT 3.970 15.410 4.410 16.560 ;
        RECT 10.720 15.410 11.160 16.560 ;
        RECT 3.970 14.760 5.120 15.410 ;
        RECT 10.010 14.760 11.160 15.410 ;
        RECT 3.970 13.610 4.410 14.760 ;
        RECT 10.720 13.610 11.160 14.760 ;
        RECT 3.970 13.510 4.420 13.610 ;
        RECT 3.270 13.430 4.420 13.510 ;
        RECT 10.710 13.510 11.160 13.610 ;
        RECT 17.470 16.560 17.920 16.660 ;
        RECT 24.210 16.660 25.360 16.740 ;
        RECT 30.270 16.960 30.720 17.110 ;
        RECT 30.970 17.000 31.420 17.110 ;
        RECT 31.670 17.000 32.080 17.100 ;
        RECT 30.970 16.960 32.080 17.000 ;
        RECT 30.270 16.740 32.080 16.960 ;
        RECT 30.270 16.660 31.420 16.740 ;
        RECT 31.670 16.680 32.080 16.740 ;
        RECT 37.050 17.000 37.460 17.100 ;
        RECT 37.710 17.000 38.160 17.110 ;
        RECT 37.050 16.960 38.160 17.000 ;
        RECT 38.410 16.960 38.860 17.110 ;
        RECT 37.050 16.740 38.860 16.960 ;
        RECT 37.050 16.680 37.460 16.740 ;
        RECT 24.210 16.560 24.660 16.660 ;
        RECT 17.470 15.410 17.910 16.560 ;
        RECT 24.220 15.410 24.660 16.560 ;
        RECT 17.470 14.760 18.620 15.410 ;
        RECT 23.510 14.760 24.660 15.410 ;
        RECT 17.470 13.610 17.910 14.760 ;
        RECT 24.220 13.610 24.660 14.760 ;
        RECT 17.470 13.510 17.920 13.610 ;
        RECT 4.670 13.430 5.080 13.490 ;
        RECT 3.270 13.130 5.080 13.430 ;
        RECT 3.270 13.050 4.420 13.130 ;
        RECT 4.670 13.070 5.080 13.130 ;
        RECT 10.050 13.430 10.460 13.490 ;
        RECT 10.710 13.430 11.860 13.510 ;
        RECT 10.050 13.130 11.860 13.430 ;
        RECT 10.050 13.070 10.460 13.130 ;
        RECT 3.970 12.950 4.420 13.050 ;
        RECT 10.710 13.050 11.860 13.130 ;
        RECT 16.770 13.430 17.920 13.510 ;
        RECT 24.210 13.510 24.660 13.610 ;
        RECT 30.970 16.560 31.420 16.660 ;
        RECT 37.710 16.660 38.860 16.740 ;
        RECT 43.770 16.960 44.220 17.110 ;
        RECT 44.470 17.000 44.920 17.110 ;
        RECT 45.170 17.000 45.580 17.100 ;
        RECT 44.470 16.960 45.580 17.000 ;
        RECT 43.770 16.740 45.580 16.960 ;
        RECT 43.770 16.660 44.920 16.740 ;
        RECT 45.170 16.680 45.580 16.740 ;
        RECT 50.550 17.000 50.960 17.100 ;
        RECT 51.210 17.000 51.660 17.110 ;
        RECT 50.550 16.960 51.660 17.000 ;
        RECT 51.910 16.960 52.360 17.110 ;
        RECT 50.550 16.740 52.360 16.960 ;
        RECT 50.550 16.680 50.960 16.740 ;
        RECT 37.710 16.560 38.160 16.660 ;
        RECT 30.970 15.410 31.410 16.560 ;
        RECT 37.720 15.410 38.160 16.560 ;
        RECT 30.970 14.760 32.120 15.410 ;
        RECT 37.010 14.760 38.160 15.410 ;
        RECT 30.970 13.610 31.410 14.760 ;
        RECT 37.720 13.610 38.160 14.760 ;
        RECT 30.970 13.510 31.420 13.610 ;
        RECT 18.170 13.430 18.580 13.490 ;
        RECT 16.770 13.130 18.580 13.430 ;
        RECT 16.770 13.050 17.920 13.130 ;
        RECT 18.170 13.070 18.580 13.130 ;
        RECT 23.550 13.430 23.960 13.490 ;
        RECT 24.210 13.430 25.360 13.510 ;
        RECT 23.550 13.130 25.360 13.430 ;
        RECT 23.550 13.070 23.960 13.130 ;
        RECT 10.710 12.950 11.160 13.050 ;
        RECT 3.970 11.800 4.410 12.950 ;
        RECT 10.720 11.800 11.160 12.950 ;
        RECT 3.970 11.150 5.120 11.800 ;
        RECT 10.010 11.150 11.160 11.800 ;
        RECT 3.970 10.000 4.410 11.150 ;
        RECT 10.720 10.000 11.160 11.150 ;
        RECT 3.970 9.900 4.420 10.000 ;
        RECT 3.270 9.820 4.420 9.900 ;
        RECT 10.710 9.900 11.160 10.000 ;
        RECT 17.470 12.950 17.920 13.050 ;
        RECT 24.210 13.050 25.360 13.130 ;
        RECT 30.270 13.430 31.420 13.510 ;
        RECT 37.710 13.510 38.160 13.610 ;
        RECT 44.470 16.560 44.920 16.660 ;
        RECT 51.210 16.660 52.360 16.740 ;
        RECT 57.270 16.960 57.720 17.110 ;
        RECT 57.970 17.000 58.420 17.110 ;
        RECT 58.670 17.000 59.080 17.100 ;
        RECT 57.970 16.960 59.080 17.000 ;
        RECT 57.270 16.740 59.080 16.960 ;
        RECT 57.270 16.660 58.420 16.740 ;
        RECT 58.670 16.680 59.080 16.740 ;
        RECT 64.050 17.000 64.460 17.100 ;
        RECT 64.710 17.000 65.160 17.110 ;
        RECT 64.050 16.960 65.160 17.000 ;
        RECT 65.410 16.960 65.860 17.110 ;
        RECT 64.050 16.740 65.860 16.960 ;
        RECT 64.050 16.680 64.460 16.740 ;
        RECT 51.210 16.560 51.660 16.660 ;
        RECT 44.470 15.410 44.910 16.560 ;
        RECT 51.220 15.410 51.660 16.560 ;
        RECT 44.470 14.760 45.620 15.410 ;
        RECT 50.510 14.760 51.660 15.410 ;
        RECT 44.470 13.610 44.910 14.760 ;
        RECT 51.220 13.610 51.660 14.760 ;
        RECT 44.470 13.510 44.920 13.610 ;
        RECT 31.670 13.430 32.080 13.490 ;
        RECT 30.270 13.130 32.080 13.430 ;
        RECT 30.270 13.050 31.420 13.130 ;
        RECT 31.670 13.070 32.080 13.130 ;
        RECT 37.050 13.430 37.460 13.490 ;
        RECT 37.710 13.430 38.860 13.510 ;
        RECT 37.050 13.130 38.860 13.430 ;
        RECT 37.050 13.070 37.460 13.130 ;
        RECT 24.210 12.950 24.660 13.050 ;
        RECT 17.470 11.800 17.910 12.950 ;
        RECT 24.220 11.800 24.660 12.950 ;
        RECT 17.470 11.150 18.620 11.800 ;
        RECT 23.510 11.150 24.660 11.800 ;
        RECT 17.470 10.000 17.910 11.150 ;
        RECT 24.220 10.000 24.660 11.150 ;
        RECT 17.470 9.900 17.920 10.000 ;
        RECT 4.670 9.820 5.080 9.880 ;
        RECT 3.270 9.520 5.080 9.820 ;
        RECT 3.270 9.440 4.420 9.520 ;
        RECT 4.670 9.460 5.080 9.520 ;
        RECT 10.050 9.820 10.460 9.880 ;
        RECT 10.710 9.820 11.860 9.900 ;
        RECT 10.050 9.520 11.860 9.820 ;
        RECT 10.050 9.460 10.460 9.520 ;
        RECT 3.970 9.340 4.420 9.440 ;
        RECT 10.710 9.440 11.860 9.520 ;
        RECT 16.770 9.820 17.920 9.900 ;
        RECT 24.210 9.900 24.660 10.000 ;
        RECT 30.970 12.950 31.420 13.050 ;
        RECT 37.710 13.050 38.860 13.130 ;
        RECT 43.770 13.430 44.920 13.510 ;
        RECT 51.210 13.510 51.660 13.610 ;
        RECT 57.970 16.560 58.420 16.660 ;
        RECT 64.710 16.660 65.860 16.740 ;
        RECT 70.770 16.960 71.220 17.110 ;
        RECT 71.470 17.000 71.920 17.110 ;
        RECT 72.170 17.000 72.580 17.100 ;
        RECT 71.470 16.960 72.580 17.000 ;
        RECT 70.770 16.740 72.580 16.960 ;
        RECT 70.770 16.660 71.920 16.740 ;
        RECT 72.170 16.680 72.580 16.740 ;
        RECT 77.550 17.000 77.960 17.100 ;
        RECT 78.210 17.000 78.660 17.110 ;
        RECT 77.550 16.960 78.660 17.000 ;
        RECT 78.910 16.960 79.360 17.110 ;
        RECT 77.550 16.740 79.360 16.960 ;
        RECT 77.550 16.680 77.960 16.740 ;
        RECT 64.710 16.560 65.160 16.660 ;
        RECT 57.970 15.410 58.410 16.560 ;
        RECT 64.720 15.410 65.160 16.560 ;
        RECT 57.970 14.760 59.120 15.410 ;
        RECT 64.010 14.760 65.160 15.410 ;
        RECT 57.970 13.610 58.410 14.760 ;
        RECT 64.720 13.610 65.160 14.760 ;
        RECT 57.970 13.510 58.420 13.610 ;
        RECT 45.170 13.430 45.580 13.490 ;
        RECT 43.770 13.130 45.580 13.430 ;
        RECT 43.770 13.050 44.920 13.130 ;
        RECT 45.170 13.070 45.580 13.130 ;
        RECT 50.550 13.430 50.960 13.490 ;
        RECT 51.210 13.430 52.360 13.510 ;
        RECT 50.550 13.130 52.360 13.430 ;
        RECT 50.550 13.070 50.960 13.130 ;
        RECT 37.710 12.950 38.160 13.050 ;
        RECT 30.970 11.800 31.410 12.950 ;
        RECT 37.720 11.800 38.160 12.950 ;
        RECT 30.970 11.150 32.120 11.800 ;
        RECT 37.010 11.150 38.160 11.800 ;
        RECT 30.970 10.000 31.410 11.150 ;
        RECT 37.720 10.000 38.160 11.150 ;
        RECT 30.970 9.900 31.420 10.000 ;
        RECT 18.170 9.820 18.580 9.880 ;
        RECT 16.770 9.520 18.580 9.820 ;
        RECT 16.770 9.440 17.920 9.520 ;
        RECT 18.170 9.460 18.580 9.520 ;
        RECT 23.550 9.820 23.960 9.880 ;
        RECT 24.210 9.820 25.360 9.900 ;
        RECT 23.550 9.520 25.360 9.820 ;
        RECT 23.550 9.460 23.960 9.520 ;
        RECT 10.710 9.340 11.160 9.440 ;
        RECT 3.970 8.190 4.410 9.340 ;
        RECT 10.720 8.190 11.160 9.340 ;
        RECT 3.970 7.540 5.120 8.190 ;
        RECT 10.010 7.540 11.160 8.190 ;
        RECT 3.970 6.390 4.410 7.540 ;
        RECT 10.720 6.390 11.160 7.540 ;
        RECT 3.970 6.290 4.420 6.390 ;
        RECT 3.270 6.210 4.420 6.290 ;
        RECT 10.710 6.290 11.160 6.390 ;
        RECT 17.470 9.340 17.920 9.440 ;
        RECT 24.210 9.440 25.360 9.520 ;
        RECT 30.270 9.820 31.420 9.900 ;
        RECT 37.710 9.900 38.160 10.000 ;
        RECT 44.470 12.950 44.920 13.050 ;
        RECT 51.210 13.050 52.360 13.130 ;
        RECT 57.270 13.430 58.420 13.510 ;
        RECT 64.710 13.510 65.160 13.610 ;
        RECT 71.470 16.560 71.920 16.660 ;
        RECT 78.210 16.660 79.360 16.740 ;
        RECT 84.270 16.960 84.720 17.110 ;
        RECT 84.970 17.000 85.420 17.110 ;
        RECT 85.670 17.000 86.080 17.100 ;
        RECT 84.970 16.960 86.080 17.000 ;
        RECT 84.270 16.740 86.080 16.960 ;
        RECT 84.270 16.660 85.420 16.740 ;
        RECT 85.670 16.680 86.080 16.740 ;
        RECT 91.050 17.000 91.460 17.100 ;
        RECT 91.710 17.000 92.160 17.110 ;
        RECT 91.050 16.960 92.160 17.000 ;
        RECT 92.410 16.960 92.860 17.110 ;
        RECT 91.050 16.740 92.860 16.960 ;
        RECT 91.050 16.680 91.460 16.740 ;
        RECT 78.210 16.560 78.660 16.660 ;
        RECT 71.470 15.410 71.910 16.560 ;
        RECT 78.220 15.410 78.660 16.560 ;
        RECT 71.470 14.760 72.620 15.410 ;
        RECT 77.510 14.760 78.660 15.410 ;
        RECT 71.470 13.610 71.910 14.760 ;
        RECT 78.220 13.610 78.660 14.760 ;
        RECT 71.470 13.510 71.920 13.610 ;
        RECT 58.670 13.430 59.080 13.490 ;
        RECT 57.270 13.130 59.080 13.430 ;
        RECT 57.270 13.050 58.420 13.130 ;
        RECT 58.670 13.070 59.080 13.130 ;
        RECT 64.050 13.430 64.460 13.490 ;
        RECT 64.710 13.430 65.860 13.510 ;
        RECT 64.050 13.130 65.860 13.430 ;
        RECT 64.050 13.070 64.460 13.130 ;
        RECT 51.210 12.950 51.660 13.050 ;
        RECT 44.470 11.800 44.910 12.950 ;
        RECT 51.220 11.800 51.660 12.950 ;
        RECT 44.470 11.150 45.620 11.800 ;
        RECT 50.510 11.150 51.660 11.800 ;
        RECT 44.470 10.000 44.910 11.150 ;
        RECT 51.220 10.000 51.660 11.150 ;
        RECT 44.470 9.900 44.920 10.000 ;
        RECT 31.670 9.820 32.080 9.880 ;
        RECT 30.270 9.520 32.080 9.820 ;
        RECT 30.270 9.440 31.420 9.520 ;
        RECT 31.670 9.460 32.080 9.520 ;
        RECT 37.050 9.820 37.460 9.880 ;
        RECT 37.710 9.820 38.860 9.900 ;
        RECT 37.050 9.520 38.860 9.820 ;
        RECT 37.050 9.460 37.460 9.520 ;
        RECT 24.210 9.340 24.660 9.440 ;
        RECT 17.470 8.190 17.910 9.340 ;
        RECT 24.220 8.190 24.660 9.340 ;
        RECT 17.470 7.540 18.620 8.190 ;
        RECT 23.510 7.540 24.660 8.190 ;
        RECT 17.470 6.390 17.910 7.540 ;
        RECT 24.220 6.390 24.660 7.540 ;
        RECT 17.470 6.290 17.920 6.390 ;
        RECT 4.670 6.210 5.080 6.270 ;
        RECT 3.270 5.910 5.080 6.210 ;
        RECT 3.270 5.830 4.420 5.910 ;
        RECT 4.670 5.850 5.080 5.910 ;
        RECT 10.050 6.210 10.460 6.270 ;
        RECT 10.710 6.210 11.860 6.290 ;
        RECT 10.050 5.910 11.860 6.210 ;
        RECT 10.050 5.850 10.460 5.910 ;
        RECT 3.970 5.730 4.420 5.830 ;
        RECT 10.710 5.830 11.860 5.910 ;
        RECT 16.770 6.210 17.920 6.290 ;
        RECT 24.210 6.290 24.660 6.390 ;
        RECT 30.970 9.340 31.420 9.440 ;
        RECT 37.710 9.440 38.860 9.520 ;
        RECT 43.770 9.820 44.920 9.900 ;
        RECT 51.210 9.900 51.660 10.000 ;
        RECT 57.970 12.950 58.420 13.050 ;
        RECT 64.710 13.050 65.860 13.130 ;
        RECT 70.770 13.430 71.920 13.510 ;
        RECT 78.210 13.510 78.660 13.610 ;
        RECT 84.970 16.560 85.420 16.660 ;
        RECT 91.710 16.660 92.860 16.740 ;
        RECT 97.770 16.960 98.220 17.110 ;
        RECT 98.470 17.000 98.920 17.110 ;
        RECT 99.170 17.000 99.580 17.100 ;
        RECT 98.470 16.960 99.580 17.000 ;
        RECT 97.770 16.740 99.580 16.960 ;
        RECT 97.770 16.660 98.920 16.740 ;
        RECT 99.170 16.680 99.580 16.740 ;
        RECT 104.550 17.000 104.960 17.100 ;
        RECT 105.210 17.000 105.660 17.110 ;
        RECT 104.550 16.960 105.660 17.000 ;
        RECT 105.910 16.960 106.360 17.110 ;
        RECT 104.550 16.740 106.360 16.960 ;
        RECT 104.550 16.680 104.960 16.740 ;
        RECT 91.710 16.560 92.160 16.660 ;
        RECT 84.970 15.410 85.410 16.560 ;
        RECT 91.720 15.410 92.160 16.560 ;
        RECT 84.970 14.760 86.120 15.410 ;
        RECT 91.010 14.760 92.160 15.410 ;
        RECT 84.970 13.610 85.410 14.760 ;
        RECT 91.720 13.610 92.160 14.760 ;
        RECT 84.970 13.510 85.420 13.610 ;
        RECT 72.170 13.430 72.580 13.490 ;
        RECT 70.770 13.130 72.580 13.430 ;
        RECT 70.770 13.050 71.920 13.130 ;
        RECT 72.170 13.070 72.580 13.130 ;
        RECT 77.550 13.430 77.960 13.490 ;
        RECT 78.210 13.430 79.360 13.510 ;
        RECT 77.550 13.130 79.360 13.430 ;
        RECT 77.550 13.070 77.960 13.130 ;
        RECT 64.710 12.950 65.160 13.050 ;
        RECT 57.970 11.800 58.410 12.950 ;
        RECT 64.720 11.800 65.160 12.950 ;
        RECT 57.970 11.150 59.120 11.800 ;
        RECT 64.010 11.150 65.160 11.800 ;
        RECT 57.970 10.000 58.410 11.150 ;
        RECT 64.720 10.000 65.160 11.150 ;
        RECT 57.970 9.900 58.420 10.000 ;
        RECT 45.170 9.820 45.580 9.880 ;
        RECT 43.770 9.520 45.580 9.820 ;
        RECT 43.770 9.440 44.920 9.520 ;
        RECT 45.170 9.460 45.580 9.520 ;
        RECT 50.550 9.820 50.960 9.880 ;
        RECT 51.210 9.820 52.360 9.900 ;
        RECT 50.550 9.520 52.360 9.820 ;
        RECT 50.550 9.460 50.960 9.520 ;
        RECT 37.710 9.340 38.160 9.440 ;
        RECT 30.970 8.190 31.410 9.340 ;
        RECT 37.720 8.190 38.160 9.340 ;
        RECT 30.970 7.540 32.120 8.190 ;
        RECT 37.010 7.540 38.160 8.190 ;
        RECT 30.970 6.390 31.410 7.540 ;
        RECT 37.720 6.390 38.160 7.540 ;
        RECT 30.970 6.290 31.420 6.390 ;
        RECT 18.170 6.210 18.580 6.270 ;
        RECT 16.770 5.910 18.580 6.210 ;
        RECT 16.770 5.830 17.920 5.910 ;
        RECT 18.170 5.850 18.580 5.910 ;
        RECT 23.550 6.210 23.960 6.270 ;
        RECT 24.210 6.210 25.360 6.290 ;
        RECT 23.550 5.910 25.360 6.210 ;
        RECT 23.550 5.850 23.960 5.910 ;
        RECT 10.710 5.730 11.160 5.830 ;
        RECT 3.970 4.580 4.410 5.730 ;
        RECT 10.720 4.580 11.160 5.730 ;
        RECT 3.970 3.930 5.120 4.580 ;
        RECT 10.010 3.930 11.160 4.580 ;
        RECT 3.970 2.780 4.410 3.930 ;
        RECT 10.720 2.780 11.160 3.930 ;
        RECT 3.970 2.680 4.420 2.780 ;
        RECT 3.270 2.600 4.420 2.680 ;
        RECT 10.710 2.680 11.160 2.780 ;
        RECT 17.470 5.730 17.920 5.830 ;
        RECT 24.210 5.830 25.360 5.910 ;
        RECT 30.270 6.210 31.420 6.290 ;
        RECT 37.710 6.290 38.160 6.390 ;
        RECT 44.470 9.340 44.920 9.440 ;
        RECT 51.210 9.440 52.360 9.520 ;
        RECT 57.270 9.820 58.420 9.900 ;
        RECT 64.710 9.900 65.160 10.000 ;
        RECT 71.470 12.950 71.920 13.050 ;
        RECT 78.210 13.050 79.360 13.130 ;
        RECT 84.270 13.430 85.420 13.510 ;
        RECT 91.710 13.510 92.160 13.610 ;
        RECT 98.470 16.560 98.920 16.660 ;
        RECT 105.210 16.660 106.360 16.740 ;
        RECT 111.270 16.960 111.720 17.110 ;
        RECT 111.970 17.000 112.420 17.110 ;
        RECT 112.670 17.000 113.080 17.100 ;
        RECT 111.970 16.960 113.080 17.000 ;
        RECT 111.270 16.740 113.080 16.960 ;
        RECT 111.270 16.660 112.420 16.740 ;
        RECT 112.670 16.680 113.080 16.740 ;
        RECT 118.050 17.000 118.460 17.100 ;
        RECT 118.710 17.000 119.160 17.110 ;
        RECT 118.050 16.960 119.160 17.000 ;
        RECT 119.410 16.960 119.860 17.110 ;
        RECT 118.050 16.740 119.860 16.960 ;
        RECT 118.050 16.680 118.460 16.740 ;
        RECT 105.210 16.560 105.660 16.660 ;
        RECT 98.470 15.410 98.910 16.560 ;
        RECT 105.220 15.410 105.660 16.560 ;
        RECT 98.470 14.760 99.620 15.410 ;
        RECT 104.510 14.760 105.660 15.410 ;
        RECT 98.470 13.610 98.910 14.760 ;
        RECT 105.220 13.610 105.660 14.760 ;
        RECT 98.470 13.510 98.920 13.610 ;
        RECT 85.670 13.430 86.080 13.490 ;
        RECT 84.270 13.130 86.080 13.430 ;
        RECT 84.270 13.050 85.420 13.130 ;
        RECT 85.670 13.070 86.080 13.130 ;
        RECT 91.050 13.430 91.460 13.490 ;
        RECT 91.710 13.430 92.860 13.510 ;
        RECT 91.050 13.130 92.860 13.430 ;
        RECT 91.050 13.070 91.460 13.130 ;
        RECT 78.210 12.950 78.660 13.050 ;
        RECT 71.470 11.800 71.910 12.950 ;
        RECT 78.220 11.800 78.660 12.950 ;
        RECT 71.470 11.150 72.620 11.800 ;
        RECT 77.510 11.150 78.660 11.800 ;
        RECT 71.470 10.000 71.910 11.150 ;
        RECT 78.220 10.000 78.660 11.150 ;
        RECT 71.470 9.900 71.920 10.000 ;
        RECT 58.670 9.820 59.080 9.880 ;
        RECT 57.270 9.520 59.080 9.820 ;
        RECT 57.270 9.440 58.420 9.520 ;
        RECT 58.670 9.460 59.080 9.520 ;
        RECT 64.050 9.820 64.460 9.880 ;
        RECT 64.710 9.820 65.860 9.900 ;
        RECT 64.050 9.520 65.860 9.820 ;
        RECT 64.050 9.460 64.460 9.520 ;
        RECT 51.210 9.340 51.660 9.440 ;
        RECT 44.470 8.190 44.910 9.340 ;
        RECT 51.220 8.190 51.660 9.340 ;
        RECT 44.470 7.540 45.620 8.190 ;
        RECT 50.510 7.540 51.660 8.190 ;
        RECT 44.470 6.390 44.910 7.540 ;
        RECT 51.220 6.390 51.660 7.540 ;
        RECT 44.470 6.290 44.920 6.390 ;
        RECT 31.670 6.210 32.080 6.270 ;
        RECT 30.270 5.910 32.080 6.210 ;
        RECT 30.270 5.830 31.420 5.910 ;
        RECT 31.670 5.850 32.080 5.910 ;
        RECT 37.050 6.210 37.460 6.270 ;
        RECT 37.710 6.210 38.860 6.290 ;
        RECT 37.050 5.910 38.860 6.210 ;
        RECT 37.050 5.850 37.460 5.910 ;
        RECT 24.210 5.730 24.660 5.830 ;
        RECT 17.470 4.580 17.910 5.730 ;
        RECT 24.220 4.580 24.660 5.730 ;
        RECT 17.470 3.930 18.620 4.580 ;
        RECT 23.510 3.930 24.660 4.580 ;
        RECT 17.470 2.780 17.910 3.930 ;
        RECT 24.220 2.780 24.660 3.930 ;
        RECT 17.470 2.680 17.920 2.780 ;
        RECT 4.670 2.600 5.080 2.660 ;
        RECT 3.270 2.300 5.080 2.600 ;
        RECT 3.270 2.220 4.420 2.300 ;
        RECT 4.670 2.240 5.080 2.300 ;
        RECT 10.050 2.600 10.460 2.660 ;
        RECT 10.710 2.600 11.860 2.680 ;
        RECT 10.050 2.300 11.860 2.600 ;
        RECT 10.050 2.240 10.460 2.300 ;
        RECT 3.970 2.120 4.420 2.220 ;
        RECT 10.710 2.220 11.860 2.300 ;
        RECT 16.770 2.600 17.920 2.680 ;
        RECT 24.210 2.680 24.660 2.780 ;
        RECT 30.970 5.730 31.420 5.830 ;
        RECT 37.710 5.830 38.860 5.910 ;
        RECT 43.770 6.210 44.920 6.290 ;
        RECT 51.210 6.290 51.660 6.390 ;
        RECT 57.970 9.340 58.420 9.440 ;
        RECT 64.710 9.440 65.860 9.520 ;
        RECT 70.770 9.820 71.920 9.900 ;
        RECT 78.210 9.900 78.660 10.000 ;
        RECT 84.970 12.950 85.420 13.050 ;
        RECT 91.710 13.050 92.860 13.130 ;
        RECT 97.770 13.430 98.920 13.510 ;
        RECT 105.210 13.510 105.660 13.610 ;
        RECT 111.970 16.560 112.420 16.660 ;
        RECT 118.710 16.660 119.860 16.740 ;
        RECT 124.770 16.960 125.220 17.110 ;
        RECT 125.470 17.000 125.920 17.110 ;
        RECT 126.170 17.000 126.580 17.100 ;
        RECT 125.470 16.960 126.580 17.000 ;
        RECT 124.770 16.740 126.580 16.960 ;
        RECT 124.770 16.660 125.920 16.740 ;
        RECT 126.170 16.680 126.580 16.740 ;
        RECT 131.550 17.000 131.960 17.100 ;
        RECT 132.210 17.000 132.660 17.110 ;
        RECT 131.550 16.960 132.660 17.000 ;
        RECT 132.910 16.960 133.360 17.110 ;
        RECT 131.550 16.740 133.360 16.960 ;
        RECT 131.550 16.680 131.960 16.740 ;
        RECT 118.710 16.560 119.160 16.660 ;
        RECT 111.970 15.410 112.410 16.560 ;
        RECT 118.720 15.410 119.160 16.560 ;
        RECT 111.970 14.760 113.120 15.410 ;
        RECT 118.010 14.760 119.160 15.410 ;
        RECT 111.970 13.610 112.410 14.760 ;
        RECT 118.720 13.610 119.160 14.760 ;
        RECT 111.970 13.510 112.420 13.610 ;
        RECT 99.170 13.430 99.580 13.490 ;
        RECT 97.770 13.130 99.580 13.430 ;
        RECT 97.770 13.050 98.920 13.130 ;
        RECT 99.170 13.070 99.580 13.130 ;
        RECT 104.550 13.430 104.960 13.490 ;
        RECT 105.210 13.430 106.360 13.510 ;
        RECT 104.550 13.130 106.360 13.430 ;
        RECT 104.550 13.070 104.960 13.130 ;
        RECT 91.710 12.950 92.160 13.050 ;
        RECT 84.970 11.800 85.410 12.950 ;
        RECT 91.720 11.800 92.160 12.950 ;
        RECT 84.970 11.150 86.120 11.800 ;
        RECT 91.010 11.150 92.160 11.800 ;
        RECT 84.970 10.000 85.410 11.150 ;
        RECT 91.720 10.000 92.160 11.150 ;
        RECT 84.970 9.900 85.420 10.000 ;
        RECT 72.170 9.820 72.580 9.880 ;
        RECT 70.770 9.520 72.580 9.820 ;
        RECT 70.770 9.440 71.920 9.520 ;
        RECT 72.170 9.460 72.580 9.520 ;
        RECT 77.550 9.820 77.960 9.880 ;
        RECT 78.210 9.820 79.360 9.900 ;
        RECT 77.550 9.520 79.360 9.820 ;
        RECT 77.550 9.460 77.960 9.520 ;
        RECT 64.710 9.340 65.160 9.440 ;
        RECT 57.970 8.190 58.410 9.340 ;
        RECT 64.720 8.190 65.160 9.340 ;
        RECT 57.970 7.540 59.120 8.190 ;
        RECT 64.010 7.540 65.160 8.190 ;
        RECT 57.970 6.390 58.410 7.540 ;
        RECT 64.720 6.390 65.160 7.540 ;
        RECT 57.970 6.290 58.420 6.390 ;
        RECT 45.170 6.210 45.580 6.270 ;
        RECT 43.770 5.910 45.580 6.210 ;
        RECT 43.770 5.830 44.920 5.910 ;
        RECT 45.170 5.850 45.580 5.910 ;
        RECT 50.550 6.210 50.960 6.270 ;
        RECT 51.210 6.210 52.360 6.290 ;
        RECT 50.550 5.910 52.360 6.210 ;
        RECT 50.550 5.850 50.960 5.910 ;
        RECT 37.710 5.730 38.160 5.830 ;
        RECT 30.970 4.580 31.410 5.730 ;
        RECT 37.720 4.580 38.160 5.730 ;
        RECT 30.970 3.930 32.120 4.580 ;
        RECT 37.010 3.930 38.160 4.580 ;
        RECT 30.970 2.780 31.410 3.930 ;
        RECT 37.720 2.780 38.160 3.930 ;
        RECT 30.970 2.680 31.420 2.780 ;
        RECT 18.170 2.600 18.580 2.660 ;
        RECT 16.770 2.300 18.580 2.600 ;
        RECT 16.770 2.220 17.920 2.300 ;
        RECT 18.170 2.240 18.580 2.300 ;
        RECT 23.550 2.600 23.960 2.660 ;
        RECT 24.210 2.600 25.360 2.680 ;
        RECT 23.550 2.300 25.360 2.600 ;
        RECT 23.550 2.240 23.960 2.300 ;
        RECT 10.710 2.120 11.160 2.220 ;
        RECT 3.970 0.970 4.410 2.120 ;
        RECT 10.720 0.970 11.160 2.120 ;
        RECT 3.970 0.320 5.120 0.970 ;
        RECT 10.010 0.320 11.160 0.970 ;
        RECT 3.970 -0.830 4.410 0.320 ;
        RECT 10.720 -0.830 11.160 0.320 ;
        RECT 3.970 -0.930 4.420 -0.830 ;
        RECT 3.270 -1.010 4.420 -0.930 ;
        RECT 10.710 -0.930 11.160 -0.830 ;
        RECT 17.470 2.120 17.920 2.220 ;
        RECT 24.210 2.220 25.360 2.300 ;
        RECT 30.270 2.600 31.420 2.680 ;
        RECT 37.710 2.680 38.160 2.780 ;
        RECT 44.470 5.730 44.920 5.830 ;
        RECT 51.210 5.830 52.360 5.910 ;
        RECT 57.270 6.210 58.420 6.290 ;
        RECT 64.710 6.290 65.160 6.390 ;
        RECT 71.470 9.340 71.920 9.440 ;
        RECT 78.210 9.440 79.360 9.520 ;
        RECT 84.270 9.820 85.420 9.900 ;
        RECT 91.710 9.900 92.160 10.000 ;
        RECT 98.470 12.950 98.920 13.050 ;
        RECT 105.210 13.050 106.360 13.130 ;
        RECT 111.270 13.430 112.420 13.510 ;
        RECT 118.710 13.510 119.160 13.610 ;
        RECT 125.470 16.560 125.920 16.660 ;
        RECT 132.210 16.660 133.360 16.740 ;
        RECT 138.270 16.960 138.720 17.110 ;
        RECT 138.970 17.000 139.420 17.110 ;
        RECT 139.670 17.000 140.080 17.100 ;
        RECT 138.970 16.960 140.080 17.000 ;
        RECT 138.270 16.740 140.080 16.960 ;
        RECT 138.270 16.660 139.420 16.740 ;
        RECT 139.670 16.680 140.080 16.740 ;
        RECT 145.050 17.000 145.460 17.100 ;
        RECT 145.710 17.000 146.160 17.110 ;
        RECT 145.050 16.960 146.160 17.000 ;
        RECT 146.410 16.960 146.860 17.110 ;
        RECT 145.050 16.740 146.860 16.960 ;
        RECT 145.050 16.680 145.460 16.740 ;
        RECT 132.210 16.560 132.660 16.660 ;
        RECT 125.470 15.410 125.910 16.560 ;
        RECT 132.220 15.410 132.660 16.560 ;
        RECT 125.470 14.760 126.620 15.410 ;
        RECT 131.510 14.760 132.660 15.410 ;
        RECT 125.470 13.610 125.910 14.760 ;
        RECT 132.220 13.610 132.660 14.760 ;
        RECT 125.470 13.510 125.920 13.610 ;
        RECT 112.670 13.430 113.080 13.490 ;
        RECT 111.270 13.130 113.080 13.430 ;
        RECT 111.270 13.050 112.420 13.130 ;
        RECT 112.670 13.070 113.080 13.130 ;
        RECT 118.050 13.430 118.460 13.490 ;
        RECT 118.710 13.430 119.860 13.510 ;
        RECT 118.050 13.130 119.860 13.430 ;
        RECT 118.050 13.070 118.460 13.130 ;
        RECT 105.210 12.950 105.660 13.050 ;
        RECT 98.470 11.800 98.910 12.950 ;
        RECT 105.220 11.800 105.660 12.950 ;
        RECT 98.470 11.150 99.620 11.800 ;
        RECT 104.510 11.150 105.660 11.800 ;
        RECT 98.470 10.000 98.910 11.150 ;
        RECT 105.220 10.000 105.660 11.150 ;
        RECT 98.470 9.900 98.920 10.000 ;
        RECT 85.670 9.820 86.080 9.880 ;
        RECT 84.270 9.520 86.080 9.820 ;
        RECT 84.270 9.440 85.420 9.520 ;
        RECT 85.670 9.460 86.080 9.520 ;
        RECT 91.050 9.820 91.460 9.880 ;
        RECT 91.710 9.820 92.860 9.900 ;
        RECT 91.050 9.520 92.860 9.820 ;
        RECT 91.050 9.460 91.460 9.520 ;
        RECT 78.210 9.340 78.660 9.440 ;
        RECT 71.470 8.190 71.910 9.340 ;
        RECT 78.220 8.190 78.660 9.340 ;
        RECT 71.470 7.540 72.620 8.190 ;
        RECT 77.510 7.540 78.660 8.190 ;
        RECT 71.470 6.390 71.910 7.540 ;
        RECT 78.220 6.390 78.660 7.540 ;
        RECT 71.470 6.290 71.920 6.390 ;
        RECT 58.670 6.210 59.080 6.270 ;
        RECT 57.270 5.910 59.080 6.210 ;
        RECT 57.270 5.830 58.420 5.910 ;
        RECT 58.670 5.850 59.080 5.910 ;
        RECT 64.050 6.210 64.460 6.270 ;
        RECT 64.710 6.210 65.860 6.290 ;
        RECT 64.050 5.910 65.860 6.210 ;
        RECT 64.050 5.850 64.460 5.910 ;
        RECT 51.210 5.730 51.660 5.830 ;
        RECT 44.470 4.580 44.910 5.730 ;
        RECT 51.220 4.580 51.660 5.730 ;
        RECT 44.470 3.930 45.620 4.580 ;
        RECT 50.510 3.930 51.660 4.580 ;
        RECT 44.470 2.780 44.910 3.930 ;
        RECT 51.220 2.780 51.660 3.930 ;
        RECT 44.470 2.680 44.920 2.780 ;
        RECT 31.670 2.600 32.080 2.660 ;
        RECT 30.270 2.300 32.080 2.600 ;
        RECT 30.270 2.220 31.420 2.300 ;
        RECT 31.670 2.240 32.080 2.300 ;
        RECT 37.050 2.600 37.460 2.660 ;
        RECT 37.710 2.600 38.860 2.680 ;
        RECT 37.050 2.300 38.860 2.600 ;
        RECT 37.050 2.240 37.460 2.300 ;
        RECT 24.210 2.120 24.660 2.220 ;
        RECT 17.470 0.970 17.910 2.120 ;
        RECT 24.220 0.970 24.660 2.120 ;
        RECT 17.470 0.320 18.620 0.970 ;
        RECT 23.510 0.320 24.660 0.970 ;
        RECT 17.470 -0.830 17.910 0.320 ;
        RECT 24.220 -0.830 24.660 0.320 ;
        RECT 17.470 -0.930 17.920 -0.830 ;
        RECT 4.670 -1.010 5.080 -0.950 ;
        RECT 3.270 -1.310 5.080 -1.010 ;
        RECT 3.270 -1.390 4.420 -1.310 ;
        RECT 4.670 -1.370 5.080 -1.310 ;
        RECT 10.050 -1.010 10.460 -0.950 ;
        RECT 10.710 -1.010 11.860 -0.930 ;
        RECT 10.050 -1.310 11.860 -1.010 ;
        RECT 10.050 -1.370 10.460 -1.310 ;
        RECT 3.970 -1.490 4.420 -1.390 ;
        RECT 10.710 -1.390 11.860 -1.310 ;
        RECT 16.770 -1.010 17.920 -0.930 ;
        RECT 24.210 -0.930 24.660 -0.830 ;
        RECT 30.970 2.120 31.420 2.220 ;
        RECT 37.710 2.220 38.860 2.300 ;
        RECT 43.770 2.600 44.920 2.680 ;
        RECT 51.210 2.680 51.660 2.780 ;
        RECT 57.970 5.730 58.420 5.830 ;
        RECT 64.710 5.830 65.860 5.910 ;
        RECT 70.770 6.210 71.920 6.290 ;
        RECT 78.210 6.290 78.660 6.390 ;
        RECT 84.970 9.340 85.420 9.440 ;
        RECT 91.710 9.440 92.860 9.520 ;
        RECT 97.770 9.820 98.920 9.900 ;
        RECT 105.210 9.900 105.660 10.000 ;
        RECT 111.970 12.950 112.420 13.050 ;
        RECT 118.710 13.050 119.860 13.130 ;
        RECT 124.770 13.430 125.920 13.510 ;
        RECT 132.210 13.510 132.660 13.610 ;
        RECT 138.970 16.560 139.420 16.660 ;
        RECT 145.710 16.660 146.860 16.740 ;
        RECT 151.770 16.960 152.220 17.110 ;
        RECT 152.470 17.000 152.920 17.110 ;
        RECT 153.170 17.000 153.580 17.100 ;
        RECT 152.470 16.960 153.580 17.000 ;
        RECT 151.770 16.740 153.580 16.960 ;
        RECT 151.770 16.660 152.920 16.740 ;
        RECT 153.170 16.680 153.580 16.740 ;
        RECT 158.550 17.000 158.960 17.100 ;
        RECT 159.210 17.000 159.660 17.110 ;
        RECT 158.550 16.960 159.660 17.000 ;
        RECT 159.910 16.960 160.360 17.110 ;
        RECT 158.550 16.740 160.360 16.960 ;
        RECT 158.550 16.680 158.960 16.740 ;
        RECT 145.710 16.560 146.160 16.660 ;
        RECT 138.970 15.410 139.410 16.560 ;
        RECT 145.720 15.410 146.160 16.560 ;
        RECT 138.970 14.760 140.120 15.410 ;
        RECT 145.010 14.760 146.160 15.410 ;
        RECT 138.970 13.610 139.410 14.760 ;
        RECT 145.720 13.610 146.160 14.760 ;
        RECT 138.970 13.510 139.420 13.610 ;
        RECT 126.170 13.430 126.580 13.490 ;
        RECT 124.770 13.130 126.580 13.430 ;
        RECT 124.770 13.050 125.920 13.130 ;
        RECT 126.170 13.070 126.580 13.130 ;
        RECT 131.550 13.430 131.960 13.490 ;
        RECT 132.210 13.430 133.360 13.510 ;
        RECT 131.550 13.130 133.360 13.430 ;
        RECT 131.550 13.070 131.960 13.130 ;
        RECT 118.710 12.950 119.160 13.050 ;
        RECT 111.970 11.800 112.410 12.950 ;
        RECT 118.720 11.800 119.160 12.950 ;
        RECT 111.970 11.150 113.120 11.800 ;
        RECT 118.010 11.150 119.160 11.800 ;
        RECT 111.970 10.000 112.410 11.150 ;
        RECT 118.720 10.000 119.160 11.150 ;
        RECT 111.970 9.900 112.420 10.000 ;
        RECT 99.170 9.820 99.580 9.880 ;
        RECT 97.770 9.520 99.580 9.820 ;
        RECT 97.770 9.440 98.920 9.520 ;
        RECT 99.170 9.460 99.580 9.520 ;
        RECT 104.550 9.820 104.960 9.880 ;
        RECT 105.210 9.820 106.360 9.900 ;
        RECT 104.550 9.520 106.360 9.820 ;
        RECT 104.550 9.460 104.960 9.520 ;
        RECT 91.710 9.340 92.160 9.440 ;
        RECT 84.970 8.190 85.410 9.340 ;
        RECT 91.720 8.190 92.160 9.340 ;
        RECT 84.970 7.540 86.120 8.190 ;
        RECT 91.010 7.540 92.160 8.190 ;
        RECT 84.970 6.390 85.410 7.540 ;
        RECT 91.720 6.390 92.160 7.540 ;
        RECT 84.970 6.290 85.420 6.390 ;
        RECT 72.170 6.210 72.580 6.270 ;
        RECT 70.770 5.910 72.580 6.210 ;
        RECT 70.770 5.830 71.920 5.910 ;
        RECT 72.170 5.850 72.580 5.910 ;
        RECT 77.550 6.210 77.960 6.270 ;
        RECT 78.210 6.210 79.360 6.290 ;
        RECT 77.550 5.910 79.360 6.210 ;
        RECT 77.550 5.850 77.960 5.910 ;
        RECT 64.710 5.730 65.160 5.830 ;
        RECT 57.970 4.580 58.410 5.730 ;
        RECT 64.720 4.580 65.160 5.730 ;
        RECT 57.970 3.930 59.120 4.580 ;
        RECT 64.010 3.930 65.160 4.580 ;
        RECT 57.970 2.780 58.410 3.930 ;
        RECT 64.720 2.780 65.160 3.930 ;
        RECT 57.970 2.680 58.420 2.780 ;
        RECT 45.170 2.600 45.580 2.660 ;
        RECT 43.770 2.300 45.580 2.600 ;
        RECT 43.770 2.220 44.920 2.300 ;
        RECT 45.170 2.240 45.580 2.300 ;
        RECT 50.550 2.600 50.960 2.660 ;
        RECT 51.210 2.600 52.360 2.680 ;
        RECT 50.550 2.300 52.360 2.600 ;
        RECT 50.550 2.240 50.960 2.300 ;
        RECT 37.710 2.120 38.160 2.220 ;
        RECT 30.970 0.970 31.410 2.120 ;
        RECT 37.720 0.970 38.160 2.120 ;
        RECT 30.970 0.320 32.120 0.970 ;
        RECT 37.010 0.320 38.160 0.970 ;
        RECT 30.970 -0.830 31.410 0.320 ;
        RECT 37.720 -0.830 38.160 0.320 ;
        RECT 30.970 -0.930 31.420 -0.830 ;
        RECT 18.170 -1.010 18.580 -0.950 ;
        RECT 16.770 -1.310 18.580 -1.010 ;
        RECT 16.770 -1.390 17.920 -1.310 ;
        RECT 18.170 -1.370 18.580 -1.310 ;
        RECT 23.550 -1.010 23.960 -0.950 ;
        RECT 24.210 -1.010 25.360 -0.930 ;
        RECT 23.550 -1.310 25.360 -1.010 ;
        RECT 23.550 -1.370 23.960 -1.310 ;
        RECT 10.710 -1.490 11.160 -1.390 ;
        RECT 3.970 -2.640 4.410 -1.490 ;
        RECT 10.720 -2.640 11.160 -1.490 ;
        RECT 3.970 -3.290 5.120 -2.640 ;
        RECT 10.010 -3.290 11.160 -2.640 ;
        RECT 3.970 -4.440 4.410 -3.290 ;
        RECT 10.720 -4.440 11.160 -3.290 ;
        RECT 3.970 -4.540 4.420 -4.440 ;
        RECT 3.270 -4.620 4.420 -4.540 ;
        RECT 10.710 -4.540 11.160 -4.440 ;
        RECT 17.470 -1.490 17.920 -1.390 ;
        RECT 24.210 -1.390 25.360 -1.310 ;
        RECT 30.270 -1.010 31.420 -0.930 ;
        RECT 37.710 -0.930 38.160 -0.830 ;
        RECT 44.470 2.120 44.920 2.220 ;
        RECT 51.210 2.220 52.360 2.300 ;
        RECT 57.270 2.600 58.420 2.680 ;
        RECT 64.710 2.680 65.160 2.780 ;
        RECT 71.470 5.730 71.920 5.830 ;
        RECT 78.210 5.830 79.360 5.910 ;
        RECT 84.270 6.210 85.420 6.290 ;
        RECT 91.710 6.290 92.160 6.390 ;
        RECT 98.470 9.340 98.920 9.440 ;
        RECT 105.210 9.440 106.360 9.520 ;
        RECT 111.270 9.820 112.420 9.900 ;
        RECT 118.710 9.900 119.160 10.000 ;
        RECT 125.470 12.950 125.920 13.050 ;
        RECT 132.210 13.050 133.360 13.130 ;
        RECT 138.270 13.430 139.420 13.510 ;
        RECT 145.710 13.510 146.160 13.610 ;
        RECT 152.470 16.560 152.920 16.660 ;
        RECT 159.210 16.660 160.360 16.740 ;
        RECT 165.270 16.960 165.720 17.110 ;
        RECT 165.970 17.000 166.420 17.110 ;
        RECT 166.670 17.000 167.080 17.100 ;
        RECT 165.970 16.960 167.080 17.000 ;
        RECT 165.270 16.740 167.080 16.960 ;
        RECT 165.270 16.660 166.420 16.740 ;
        RECT 166.670 16.680 167.080 16.740 ;
        RECT 172.050 17.000 172.460 17.100 ;
        RECT 172.710 17.000 173.160 17.110 ;
        RECT 172.050 16.960 173.160 17.000 ;
        RECT 173.410 16.960 173.860 17.110 ;
        RECT 172.050 16.740 173.860 16.960 ;
        RECT 172.050 16.680 172.460 16.740 ;
        RECT 159.210 16.560 159.660 16.660 ;
        RECT 152.470 15.410 152.910 16.560 ;
        RECT 159.220 15.410 159.660 16.560 ;
        RECT 152.470 14.760 153.620 15.410 ;
        RECT 158.510 14.760 159.660 15.410 ;
        RECT 152.470 13.610 152.910 14.760 ;
        RECT 159.220 13.610 159.660 14.760 ;
        RECT 152.470 13.510 152.920 13.610 ;
        RECT 139.670 13.430 140.080 13.490 ;
        RECT 138.270 13.130 140.080 13.430 ;
        RECT 138.270 13.050 139.420 13.130 ;
        RECT 139.670 13.070 140.080 13.130 ;
        RECT 145.050 13.430 145.460 13.490 ;
        RECT 145.710 13.430 146.860 13.510 ;
        RECT 145.050 13.130 146.860 13.430 ;
        RECT 145.050 13.070 145.460 13.130 ;
        RECT 132.210 12.950 132.660 13.050 ;
        RECT 125.470 11.800 125.910 12.950 ;
        RECT 132.220 11.800 132.660 12.950 ;
        RECT 125.470 11.150 126.620 11.800 ;
        RECT 131.510 11.150 132.660 11.800 ;
        RECT 125.470 10.000 125.910 11.150 ;
        RECT 132.220 10.000 132.660 11.150 ;
        RECT 125.470 9.900 125.920 10.000 ;
        RECT 112.670 9.820 113.080 9.880 ;
        RECT 111.270 9.520 113.080 9.820 ;
        RECT 111.270 9.440 112.420 9.520 ;
        RECT 112.670 9.460 113.080 9.520 ;
        RECT 118.050 9.820 118.460 9.880 ;
        RECT 118.710 9.820 119.860 9.900 ;
        RECT 118.050 9.520 119.860 9.820 ;
        RECT 118.050 9.460 118.460 9.520 ;
        RECT 105.210 9.340 105.660 9.440 ;
        RECT 98.470 8.190 98.910 9.340 ;
        RECT 105.220 8.190 105.660 9.340 ;
        RECT 98.470 7.540 99.620 8.190 ;
        RECT 104.510 7.540 105.660 8.190 ;
        RECT 98.470 6.390 98.910 7.540 ;
        RECT 105.220 6.390 105.660 7.540 ;
        RECT 98.470 6.290 98.920 6.390 ;
        RECT 85.670 6.210 86.080 6.270 ;
        RECT 84.270 5.910 86.080 6.210 ;
        RECT 84.270 5.830 85.420 5.910 ;
        RECT 85.670 5.850 86.080 5.910 ;
        RECT 91.050 6.210 91.460 6.270 ;
        RECT 91.710 6.210 92.860 6.290 ;
        RECT 91.050 5.910 92.860 6.210 ;
        RECT 91.050 5.850 91.460 5.910 ;
        RECT 78.210 5.730 78.660 5.830 ;
        RECT 71.470 4.580 71.910 5.730 ;
        RECT 78.220 4.580 78.660 5.730 ;
        RECT 71.470 3.930 72.620 4.580 ;
        RECT 77.510 3.930 78.660 4.580 ;
        RECT 71.470 2.780 71.910 3.930 ;
        RECT 78.220 2.780 78.660 3.930 ;
        RECT 71.470 2.680 71.920 2.780 ;
        RECT 58.670 2.600 59.080 2.660 ;
        RECT 57.270 2.300 59.080 2.600 ;
        RECT 57.270 2.220 58.420 2.300 ;
        RECT 58.670 2.240 59.080 2.300 ;
        RECT 64.050 2.600 64.460 2.660 ;
        RECT 64.710 2.600 65.860 2.680 ;
        RECT 64.050 2.300 65.860 2.600 ;
        RECT 64.050 2.240 64.460 2.300 ;
        RECT 51.210 2.120 51.660 2.220 ;
        RECT 44.470 0.970 44.910 2.120 ;
        RECT 51.220 0.970 51.660 2.120 ;
        RECT 44.470 0.320 45.620 0.970 ;
        RECT 50.510 0.320 51.660 0.970 ;
        RECT 44.470 -0.830 44.910 0.320 ;
        RECT 51.220 -0.830 51.660 0.320 ;
        RECT 44.470 -0.930 44.920 -0.830 ;
        RECT 31.670 -1.010 32.080 -0.950 ;
        RECT 30.270 -1.310 32.080 -1.010 ;
        RECT 30.270 -1.390 31.420 -1.310 ;
        RECT 31.670 -1.370 32.080 -1.310 ;
        RECT 37.050 -1.010 37.460 -0.950 ;
        RECT 37.710 -1.010 38.860 -0.930 ;
        RECT 37.050 -1.310 38.860 -1.010 ;
        RECT 37.050 -1.370 37.460 -1.310 ;
        RECT 24.210 -1.490 24.660 -1.390 ;
        RECT 17.470 -2.640 17.910 -1.490 ;
        RECT 24.220 -2.640 24.660 -1.490 ;
        RECT 17.470 -3.290 18.620 -2.640 ;
        RECT 23.510 -3.290 24.660 -2.640 ;
        RECT 17.470 -4.440 17.910 -3.290 ;
        RECT 24.220 -4.440 24.660 -3.290 ;
        RECT 17.470 -4.540 17.920 -4.440 ;
        RECT 4.670 -4.620 5.080 -4.560 ;
        RECT 3.270 -4.920 5.080 -4.620 ;
        RECT 3.270 -5.000 4.420 -4.920 ;
        RECT 4.670 -4.980 5.080 -4.920 ;
        RECT 10.050 -4.620 10.460 -4.560 ;
        RECT 10.710 -4.620 11.860 -4.540 ;
        RECT 10.050 -4.920 11.860 -4.620 ;
        RECT 10.050 -4.980 10.460 -4.920 ;
        RECT 3.970 -5.100 4.420 -5.000 ;
        RECT 10.710 -5.000 11.860 -4.920 ;
        RECT 16.770 -4.620 17.920 -4.540 ;
        RECT 24.210 -4.540 24.660 -4.440 ;
        RECT 30.970 -1.490 31.420 -1.390 ;
        RECT 37.710 -1.390 38.860 -1.310 ;
        RECT 43.770 -1.010 44.920 -0.930 ;
        RECT 51.210 -0.930 51.660 -0.830 ;
        RECT 57.970 2.120 58.420 2.220 ;
        RECT 64.710 2.220 65.860 2.300 ;
        RECT 70.770 2.600 71.920 2.680 ;
        RECT 78.210 2.680 78.660 2.780 ;
        RECT 84.970 5.730 85.420 5.830 ;
        RECT 91.710 5.830 92.860 5.910 ;
        RECT 97.770 6.210 98.920 6.290 ;
        RECT 105.210 6.290 105.660 6.390 ;
        RECT 111.970 9.340 112.420 9.440 ;
        RECT 118.710 9.440 119.860 9.520 ;
        RECT 124.770 9.820 125.920 9.900 ;
        RECT 132.210 9.900 132.660 10.000 ;
        RECT 138.970 12.950 139.420 13.050 ;
        RECT 145.710 13.050 146.860 13.130 ;
        RECT 151.770 13.430 152.920 13.510 ;
        RECT 159.210 13.510 159.660 13.610 ;
        RECT 165.970 16.560 166.420 16.660 ;
        RECT 172.710 16.660 173.860 16.740 ;
        RECT 178.770 16.960 179.220 17.110 ;
        RECT 179.470 17.000 179.920 17.110 ;
        RECT 180.170 17.000 180.580 17.100 ;
        RECT 179.470 16.960 180.580 17.000 ;
        RECT 178.770 16.740 180.580 16.960 ;
        RECT 178.770 16.660 179.920 16.740 ;
        RECT 180.170 16.680 180.580 16.740 ;
        RECT 185.550 17.000 185.960 17.100 ;
        RECT 186.210 17.000 186.660 17.110 ;
        RECT 185.550 16.960 186.660 17.000 ;
        RECT 186.910 16.960 187.360 17.110 ;
        RECT 185.550 16.740 187.360 16.960 ;
        RECT 185.550 16.680 185.960 16.740 ;
        RECT 172.710 16.560 173.160 16.660 ;
        RECT 165.970 15.410 166.410 16.560 ;
        RECT 172.720 15.410 173.160 16.560 ;
        RECT 165.970 14.760 167.120 15.410 ;
        RECT 172.010 14.760 173.160 15.410 ;
        RECT 165.970 13.610 166.410 14.760 ;
        RECT 172.720 13.610 173.160 14.760 ;
        RECT 165.970 13.510 166.420 13.610 ;
        RECT 153.170 13.430 153.580 13.490 ;
        RECT 151.770 13.130 153.580 13.430 ;
        RECT 151.770 13.050 152.920 13.130 ;
        RECT 153.170 13.070 153.580 13.130 ;
        RECT 158.550 13.430 158.960 13.490 ;
        RECT 159.210 13.430 160.360 13.510 ;
        RECT 158.550 13.130 160.360 13.430 ;
        RECT 158.550 13.070 158.960 13.130 ;
        RECT 145.710 12.950 146.160 13.050 ;
        RECT 138.970 11.800 139.410 12.950 ;
        RECT 145.720 11.800 146.160 12.950 ;
        RECT 138.970 11.150 140.120 11.800 ;
        RECT 145.010 11.150 146.160 11.800 ;
        RECT 138.970 10.000 139.410 11.150 ;
        RECT 145.720 10.000 146.160 11.150 ;
        RECT 138.970 9.900 139.420 10.000 ;
        RECT 126.170 9.820 126.580 9.880 ;
        RECT 124.770 9.520 126.580 9.820 ;
        RECT 124.770 9.440 125.920 9.520 ;
        RECT 126.170 9.460 126.580 9.520 ;
        RECT 131.550 9.820 131.960 9.880 ;
        RECT 132.210 9.820 133.360 9.900 ;
        RECT 131.550 9.520 133.360 9.820 ;
        RECT 131.550 9.460 131.960 9.520 ;
        RECT 118.710 9.340 119.160 9.440 ;
        RECT 111.970 8.190 112.410 9.340 ;
        RECT 118.720 8.190 119.160 9.340 ;
        RECT 111.970 7.540 113.120 8.190 ;
        RECT 118.010 7.540 119.160 8.190 ;
        RECT 111.970 6.390 112.410 7.540 ;
        RECT 118.720 6.390 119.160 7.540 ;
        RECT 111.970 6.290 112.420 6.390 ;
        RECT 99.170 6.210 99.580 6.270 ;
        RECT 97.770 5.910 99.580 6.210 ;
        RECT 97.770 5.830 98.920 5.910 ;
        RECT 99.170 5.850 99.580 5.910 ;
        RECT 104.550 6.210 104.960 6.270 ;
        RECT 105.210 6.210 106.360 6.290 ;
        RECT 104.550 5.910 106.360 6.210 ;
        RECT 104.550 5.850 104.960 5.910 ;
        RECT 91.710 5.730 92.160 5.830 ;
        RECT 84.970 4.580 85.410 5.730 ;
        RECT 91.720 4.580 92.160 5.730 ;
        RECT 84.970 3.930 86.120 4.580 ;
        RECT 91.010 3.930 92.160 4.580 ;
        RECT 84.970 2.780 85.410 3.930 ;
        RECT 91.720 2.780 92.160 3.930 ;
        RECT 84.970 2.680 85.420 2.780 ;
        RECT 72.170 2.600 72.580 2.660 ;
        RECT 70.770 2.300 72.580 2.600 ;
        RECT 70.770 2.220 71.920 2.300 ;
        RECT 72.170 2.240 72.580 2.300 ;
        RECT 77.550 2.600 77.960 2.660 ;
        RECT 78.210 2.600 79.360 2.680 ;
        RECT 77.550 2.300 79.360 2.600 ;
        RECT 77.550 2.240 77.960 2.300 ;
        RECT 64.710 2.120 65.160 2.220 ;
        RECT 57.970 0.970 58.410 2.120 ;
        RECT 64.720 0.970 65.160 2.120 ;
        RECT 57.970 0.320 59.120 0.970 ;
        RECT 64.010 0.320 65.160 0.970 ;
        RECT 57.970 -0.830 58.410 0.320 ;
        RECT 64.720 -0.830 65.160 0.320 ;
        RECT 57.970 -0.930 58.420 -0.830 ;
        RECT 45.170 -1.010 45.580 -0.950 ;
        RECT 43.770 -1.310 45.580 -1.010 ;
        RECT 43.770 -1.390 44.920 -1.310 ;
        RECT 45.170 -1.370 45.580 -1.310 ;
        RECT 50.550 -1.010 50.960 -0.950 ;
        RECT 51.210 -1.010 52.360 -0.930 ;
        RECT 50.550 -1.310 52.360 -1.010 ;
        RECT 50.550 -1.370 50.960 -1.310 ;
        RECT 37.710 -1.490 38.160 -1.390 ;
        RECT 30.970 -2.640 31.410 -1.490 ;
        RECT 37.720 -2.640 38.160 -1.490 ;
        RECT 30.970 -3.290 32.120 -2.640 ;
        RECT 37.010 -3.290 38.160 -2.640 ;
        RECT 30.970 -4.440 31.410 -3.290 ;
        RECT 37.720 -4.440 38.160 -3.290 ;
        RECT 30.970 -4.540 31.420 -4.440 ;
        RECT 18.170 -4.620 18.580 -4.560 ;
        RECT 16.770 -4.920 18.580 -4.620 ;
        RECT 16.770 -5.000 17.920 -4.920 ;
        RECT 18.170 -4.980 18.580 -4.920 ;
        RECT 23.550 -4.620 23.960 -4.560 ;
        RECT 24.210 -4.620 25.360 -4.540 ;
        RECT 23.550 -4.920 25.360 -4.620 ;
        RECT 23.550 -4.980 23.960 -4.920 ;
        RECT 10.710 -5.100 11.160 -5.000 ;
        RECT 3.970 -6.250 4.410 -5.100 ;
        RECT 10.720 -6.250 11.160 -5.100 ;
        RECT 3.970 -6.900 5.120 -6.250 ;
        RECT 10.010 -6.900 11.160 -6.250 ;
        RECT 3.970 -8.050 4.410 -6.900 ;
        RECT 10.720 -8.050 11.160 -6.900 ;
        RECT 3.970 -8.150 4.420 -8.050 ;
        RECT 3.270 -8.230 4.420 -8.150 ;
        RECT 10.710 -8.150 11.160 -8.050 ;
        RECT 17.470 -5.100 17.920 -5.000 ;
        RECT 24.210 -5.000 25.360 -4.920 ;
        RECT 30.270 -4.620 31.420 -4.540 ;
        RECT 37.710 -4.540 38.160 -4.440 ;
        RECT 44.470 -1.490 44.920 -1.390 ;
        RECT 51.210 -1.390 52.360 -1.310 ;
        RECT 57.270 -1.010 58.420 -0.930 ;
        RECT 64.710 -0.930 65.160 -0.830 ;
        RECT 71.470 2.120 71.920 2.220 ;
        RECT 78.210 2.220 79.360 2.300 ;
        RECT 84.270 2.600 85.420 2.680 ;
        RECT 91.710 2.680 92.160 2.780 ;
        RECT 98.470 5.730 98.920 5.830 ;
        RECT 105.210 5.830 106.360 5.910 ;
        RECT 111.270 6.210 112.420 6.290 ;
        RECT 118.710 6.290 119.160 6.390 ;
        RECT 125.470 9.340 125.920 9.440 ;
        RECT 132.210 9.440 133.360 9.520 ;
        RECT 138.270 9.820 139.420 9.900 ;
        RECT 145.710 9.900 146.160 10.000 ;
        RECT 152.470 12.950 152.920 13.050 ;
        RECT 159.210 13.050 160.360 13.130 ;
        RECT 165.270 13.430 166.420 13.510 ;
        RECT 172.710 13.510 173.160 13.610 ;
        RECT 179.470 16.560 179.920 16.660 ;
        RECT 186.210 16.660 187.360 16.740 ;
        RECT 192.270 16.960 192.720 17.110 ;
        RECT 192.970 17.000 193.420 17.110 ;
        RECT 193.670 17.000 194.080 17.100 ;
        RECT 192.970 16.960 194.080 17.000 ;
        RECT 192.270 16.740 194.080 16.960 ;
        RECT 192.270 16.660 193.420 16.740 ;
        RECT 193.670 16.680 194.080 16.740 ;
        RECT 199.050 17.000 199.460 17.100 ;
        RECT 199.710 17.000 200.160 17.110 ;
        RECT 199.050 16.960 200.160 17.000 ;
        RECT 200.410 16.960 200.860 17.110 ;
        RECT 199.050 16.740 200.860 16.960 ;
        RECT 199.050 16.680 199.460 16.740 ;
        RECT 186.210 16.560 186.660 16.660 ;
        RECT 179.470 15.410 179.910 16.560 ;
        RECT 186.220 15.410 186.660 16.560 ;
        RECT 179.470 14.760 180.620 15.410 ;
        RECT 185.510 14.760 186.660 15.410 ;
        RECT 179.470 13.610 179.910 14.760 ;
        RECT 186.220 13.610 186.660 14.760 ;
        RECT 179.470 13.510 179.920 13.610 ;
        RECT 166.670 13.430 167.080 13.490 ;
        RECT 165.270 13.130 167.080 13.430 ;
        RECT 165.270 13.050 166.420 13.130 ;
        RECT 166.670 13.070 167.080 13.130 ;
        RECT 172.050 13.430 172.460 13.490 ;
        RECT 172.710 13.430 173.860 13.510 ;
        RECT 172.050 13.130 173.860 13.430 ;
        RECT 172.050 13.070 172.460 13.130 ;
        RECT 159.210 12.950 159.660 13.050 ;
        RECT 152.470 11.800 152.910 12.950 ;
        RECT 159.220 11.800 159.660 12.950 ;
        RECT 152.470 11.150 153.620 11.800 ;
        RECT 158.510 11.150 159.660 11.800 ;
        RECT 152.470 10.000 152.910 11.150 ;
        RECT 159.220 10.000 159.660 11.150 ;
        RECT 152.470 9.900 152.920 10.000 ;
        RECT 139.670 9.820 140.080 9.880 ;
        RECT 138.270 9.520 140.080 9.820 ;
        RECT 138.270 9.440 139.420 9.520 ;
        RECT 139.670 9.460 140.080 9.520 ;
        RECT 145.050 9.820 145.460 9.880 ;
        RECT 145.710 9.820 146.860 9.900 ;
        RECT 145.050 9.520 146.860 9.820 ;
        RECT 145.050 9.460 145.460 9.520 ;
        RECT 132.210 9.340 132.660 9.440 ;
        RECT 125.470 8.190 125.910 9.340 ;
        RECT 132.220 8.190 132.660 9.340 ;
        RECT 125.470 7.540 126.620 8.190 ;
        RECT 131.510 7.540 132.660 8.190 ;
        RECT 125.470 6.390 125.910 7.540 ;
        RECT 132.220 6.390 132.660 7.540 ;
        RECT 125.470 6.290 125.920 6.390 ;
        RECT 112.670 6.210 113.080 6.270 ;
        RECT 111.270 5.910 113.080 6.210 ;
        RECT 111.270 5.830 112.420 5.910 ;
        RECT 112.670 5.850 113.080 5.910 ;
        RECT 118.050 6.210 118.460 6.270 ;
        RECT 118.710 6.210 119.860 6.290 ;
        RECT 118.050 5.910 119.860 6.210 ;
        RECT 118.050 5.850 118.460 5.910 ;
        RECT 105.210 5.730 105.660 5.830 ;
        RECT 98.470 4.580 98.910 5.730 ;
        RECT 105.220 4.580 105.660 5.730 ;
        RECT 98.470 3.930 99.620 4.580 ;
        RECT 104.510 3.930 105.660 4.580 ;
        RECT 98.470 2.780 98.910 3.930 ;
        RECT 105.220 2.780 105.660 3.930 ;
        RECT 98.470 2.680 98.920 2.780 ;
        RECT 85.670 2.600 86.080 2.660 ;
        RECT 84.270 2.300 86.080 2.600 ;
        RECT 84.270 2.220 85.420 2.300 ;
        RECT 85.670 2.240 86.080 2.300 ;
        RECT 91.050 2.600 91.460 2.660 ;
        RECT 91.710 2.600 92.860 2.680 ;
        RECT 91.050 2.300 92.860 2.600 ;
        RECT 91.050 2.240 91.460 2.300 ;
        RECT 78.210 2.120 78.660 2.220 ;
        RECT 71.470 0.970 71.910 2.120 ;
        RECT 78.220 0.970 78.660 2.120 ;
        RECT 71.470 0.320 72.620 0.970 ;
        RECT 77.510 0.320 78.660 0.970 ;
        RECT 71.470 -0.830 71.910 0.320 ;
        RECT 78.220 -0.830 78.660 0.320 ;
        RECT 71.470 -0.930 71.920 -0.830 ;
        RECT 58.670 -1.010 59.080 -0.950 ;
        RECT 57.270 -1.310 59.080 -1.010 ;
        RECT 57.270 -1.390 58.420 -1.310 ;
        RECT 58.670 -1.370 59.080 -1.310 ;
        RECT 64.050 -1.010 64.460 -0.950 ;
        RECT 64.710 -1.010 65.860 -0.930 ;
        RECT 64.050 -1.310 65.860 -1.010 ;
        RECT 64.050 -1.370 64.460 -1.310 ;
        RECT 51.210 -1.490 51.660 -1.390 ;
        RECT 44.470 -2.640 44.910 -1.490 ;
        RECT 51.220 -2.640 51.660 -1.490 ;
        RECT 44.470 -3.290 45.620 -2.640 ;
        RECT 50.510 -3.290 51.660 -2.640 ;
        RECT 44.470 -4.440 44.910 -3.290 ;
        RECT 51.220 -4.440 51.660 -3.290 ;
        RECT 44.470 -4.540 44.920 -4.440 ;
        RECT 31.670 -4.620 32.080 -4.560 ;
        RECT 30.270 -4.920 32.080 -4.620 ;
        RECT 30.270 -5.000 31.420 -4.920 ;
        RECT 31.670 -4.980 32.080 -4.920 ;
        RECT 37.050 -4.620 37.460 -4.560 ;
        RECT 37.710 -4.620 38.860 -4.540 ;
        RECT 37.050 -4.920 38.860 -4.620 ;
        RECT 37.050 -4.980 37.460 -4.920 ;
        RECT 24.210 -5.100 24.660 -5.000 ;
        RECT 17.470 -6.250 17.910 -5.100 ;
        RECT 24.220 -6.250 24.660 -5.100 ;
        RECT 17.470 -6.900 18.620 -6.250 ;
        RECT 23.510 -6.900 24.660 -6.250 ;
        RECT 17.470 -8.050 17.910 -6.900 ;
        RECT 24.220 -8.050 24.660 -6.900 ;
        RECT 17.470 -8.150 17.920 -8.050 ;
        RECT 4.670 -8.230 5.080 -8.170 ;
        RECT 3.270 -8.530 5.080 -8.230 ;
        RECT 3.270 -8.610 4.420 -8.530 ;
        RECT 4.670 -8.590 5.080 -8.530 ;
        RECT 10.050 -8.230 10.460 -8.170 ;
        RECT 10.710 -8.230 11.860 -8.150 ;
        RECT 10.050 -8.530 11.860 -8.230 ;
        RECT 10.050 -8.590 10.460 -8.530 ;
        RECT 3.970 -8.710 4.420 -8.610 ;
        RECT 10.710 -8.610 11.860 -8.530 ;
        RECT 16.770 -8.230 17.920 -8.150 ;
        RECT 24.210 -8.150 24.660 -8.050 ;
        RECT 30.970 -5.100 31.420 -5.000 ;
        RECT 37.710 -5.000 38.860 -4.920 ;
        RECT 43.770 -4.620 44.920 -4.540 ;
        RECT 51.210 -4.540 51.660 -4.440 ;
        RECT 57.970 -1.490 58.420 -1.390 ;
        RECT 64.710 -1.390 65.860 -1.310 ;
        RECT 70.770 -1.010 71.920 -0.930 ;
        RECT 78.210 -0.930 78.660 -0.830 ;
        RECT 84.970 2.120 85.420 2.220 ;
        RECT 91.710 2.220 92.860 2.300 ;
        RECT 97.770 2.600 98.920 2.680 ;
        RECT 105.210 2.680 105.660 2.780 ;
        RECT 111.970 5.730 112.420 5.830 ;
        RECT 118.710 5.830 119.860 5.910 ;
        RECT 124.770 6.210 125.920 6.290 ;
        RECT 132.210 6.290 132.660 6.390 ;
        RECT 138.970 9.340 139.420 9.440 ;
        RECT 145.710 9.440 146.860 9.520 ;
        RECT 151.770 9.820 152.920 9.900 ;
        RECT 159.210 9.900 159.660 10.000 ;
        RECT 165.970 12.950 166.420 13.050 ;
        RECT 172.710 13.050 173.860 13.130 ;
        RECT 178.770 13.430 179.920 13.510 ;
        RECT 186.210 13.510 186.660 13.610 ;
        RECT 192.970 16.560 193.420 16.660 ;
        RECT 199.710 16.660 200.860 16.740 ;
        RECT 205.770 16.960 206.220 17.110 ;
        RECT 206.470 17.000 206.920 17.110 ;
        RECT 207.170 17.000 207.580 17.100 ;
        RECT 206.470 16.960 207.580 17.000 ;
        RECT 205.770 16.740 207.580 16.960 ;
        RECT 205.770 16.660 206.920 16.740 ;
        RECT 207.170 16.680 207.580 16.740 ;
        RECT 212.550 17.000 212.960 17.100 ;
        RECT 213.210 17.000 213.660 17.110 ;
        RECT 212.550 16.960 213.660 17.000 ;
        RECT 213.910 16.960 214.360 17.110 ;
        RECT 212.550 16.740 214.360 16.960 ;
        RECT 212.550 16.680 212.960 16.740 ;
        RECT 199.710 16.560 200.160 16.660 ;
        RECT 192.970 15.410 193.410 16.560 ;
        RECT 199.720 15.410 200.160 16.560 ;
        RECT 192.970 14.760 194.120 15.410 ;
        RECT 199.010 14.760 200.160 15.410 ;
        RECT 192.970 13.610 193.410 14.760 ;
        RECT 199.720 13.610 200.160 14.760 ;
        RECT 192.970 13.510 193.420 13.610 ;
        RECT 180.170 13.430 180.580 13.490 ;
        RECT 178.770 13.130 180.580 13.430 ;
        RECT 178.770 13.050 179.920 13.130 ;
        RECT 180.170 13.070 180.580 13.130 ;
        RECT 185.550 13.430 185.960 13.490 ;
        RECT 186.210 13.430 187.360 13.510 ;
        RECT 185.550 13.130 187.360 13.430 ;
        RECT 185.550 13.070 185.960 13.130 ;
        RECT 172.710 12.950 173.160 13.050 ;
        RECT 165.970 11.800 166.410 12.950 ;
        RECT 172.720 11.800 173.160 12.950 ;
        RECT 165.970 11.150 167.120 11.800 ;
        RECT 172.010 11.150 173.160 11.800 ;
        RECT 165.970 10.000 166.410 11.150 ;
        RECT 172.720 10.000 173.160 11.150 ;
        RECT 165.970 9.900 166.420 10.000 ;
        RECT 153.170 9.820 153.580 9.880 ;
        RECT 151.770 9.520 153.580 9.820 ;
        RECT 151.770 9.440 152.920 9.520 ;
        RECT 153.170 9.460 153.580 9.520 ;
        RECT 158.550 9.820 158.960 9.880 ;
        RECT 159.210 9.820 160.360 9.900 ;
        RECT 158.550 9.520 160.360 9.820 ;
        RECT 158.550 9.460 158.960 9.520 ;
        RECT 145.710 9.340 146.160 9.440 ;
        RECT 138.970 8.190 139.410 9.340 ;
        RECT 145.720 8.190 146.160 9.340 ;
        RECT 138.970 7.540 140.120 8.190 ;
        RECT 145.010 7.540 146.160 8.190 ;
        RECT 138.970 6.390 139.410 7.540 ;
        RECT 145.720 6.390 146.160 7.540 ;
        RECT 138.970 6.290 139.420 6.390 ;
        RECT 126.170 6.210 126.580 6.270 ;
        RECT 124.770 5.910 126.580 6.210 ;
        RECT 124.770 5.830 125.920 5.910 ;
        RECT 126.170 5.850 126.580 5.910 ;
        RECT 131.550 6.210 131.960 6.270 ;
        RECT 132.210 6.210 133.360 6.290 ;
        RECT 131.550 5.910 133.360 6.210 ;
        RECT 131.550 5.850 131.960 5.910 ;
        RECT 118.710 5.730 119.160 5.830 ;
        RECT 111.970 4.580 112.410 5.730 ;
        RECT 118.720 4.580 119.160 5.730 ;
        RECT 111.970 3.930 113.120 4.580 ;
        RECT 118.010 3.930 119.160 4.580 ;
        RECT 111.970 2.780 112.410 3.930 ;
        RECT 118.720 2.780 119.160 3.930 ;
        RECT 111.970 2.680 112.420 2.780 ;
        RECT 99.170 2.600 99.580 2.660 ;
        RECT 97.770 2.300 99.580 2.600 ;
        RECT 97.770 2.220 98.920 2.300 ;
        RECT 99.170 2.240 99.580 2.300 ;
        RECT 104.550 2.600 104.960 2.660 ;
        RECT 105.210 2.600 106.360 2.680 ;
        RECT 104.550 2.300 106.360 2.600 ;
        RECT 104.550 2.240 104.960 2.300 ;
        RECT 91.710 2.120 92.160 2.220 ;
        RECT 84.970 0.970 85.410 2.120 ;
        RECT 91.720 0.970 92.160 2.120 ;
        RECT 84.970 0.320 86.120 0.970 ;
        RECT 91.010 0.320 92.160 0.970 ;
        RECT 84.970 -0.830 85.410 0.320 ;
        RECT 91.720 -0.830 92.160 0.320 ;
        RECT 84.970 -0.930 85.420 -0.830 ;
        RECT 72.170 -1.010 72.580 -0.950 ;
        RECT 70.770 -1.310 72.580 -1.010 ;
        RECT 70.770 -1.390 71.920 -1.310 ;
        RECT 72.170 -1.370 72.580 -1.310 ;
        RECT 77.550 -1.010 77.960 -0.950 ;
        RECT 78.210 -1.010 79.360 -0.930 ;
        RECT 77.550 -1.310 79.360 -1.010 ;
        RECT 77.550 -1.370 77.960 -1.310 ;
        RECT 64.710 -1.490 65.160 -1.390 ;
        RECT 57.970 -2.640 58.410 -1.490 ;
        RECT 64.720 -2.640 65.160 -1.490 ;
        RECT 57.970 -3.290 59.120 -2.640 ;
        RECT 64.010 -3.290 65.160 -2.640 ;
        RECT 57.970 -4.440 58.410 -3.290 ;
        RECT 64.720 -4.440 65.160 -3.290 ;
        RECT 57.970 -4.540 58.420 -4.440 ;
        RECT 45.170 -4.620 45.580 -4.560 ;
        RECT 43.770 -4.920 45.580 -4.620 ;
        RECT 43.770 -5.000 44.920 -4.920 ;
        RECT 45.170 -4.980 45.580 -4.920 ;
        RECT 50.550 -4.620 50.960 -4.560 ;
        RECT 51.210 -4.620 52.360 -4.540 ;
        RECT 50.550 -4.920 52.360 -4.620 ;
        RECT 50.550 -4.980 50.960 -4.920 ;
        RECT 37.710 -5.100 38.160 -5.000 ;
        RECT 30.970 -6.250 31.410 -5.100 ;
        RECT 37.720 -6.250 38.160 -5.100 ;
        RECT 30.970 -6.900 32.120 -6.250 ;
        RECT 37.010 -6.900 38.160 -6.250 ;
        RECT 30.970 -8.050 31.410 -6.900 ;
        RECT 37.720 -8.050 38.160 -6.900 ;
        RECT 30.970 -8.150 31.420 -8.050 ;
        RECT 18.170 -8.230 18.580 -8.170 ;
        RECT 16.770 -8.530 18.580 -8.230 ;
        RECT 16.770 -8.610 17.920 -8.530 ;
        RECT 18.170 -8.590 18.580 -8.530 ;
        RECT 23.550 -8.230 23.960 -8.170 ;
        RECT 24.210 -8.230 25.360 -8.150 ;
        RECT 23.550 -8.530 25.360 -8.230 ;
        RECT 23.550 -8.590 23.960 -8.530 ;
        RECT 10.710 -8.710 11.160 -8.610 ;
        RECT 3.970 -9.860 4.410 -8.710 ;
        RECT 10.720 -9.860 11.160 -8.710 ;
        RECT 3.970 -10.510 5.120 -9.860 ;
        RECT 10.010 -10.510 11.160 -9.860 ;
        RECT 3.970 -11.660 4.410 -10.510 ;
        RECT 10.720 -11.660 11.160 -10.510 ;
        RECT 3.970 -11.760 4.420 -11.660 ;
        RECT 3.270 -11.840 4.420 -11.760 ;
        RECT 10.710 -11.760 11.160 -11.660 ;
        RECT 17.470 -8.710 17.920 -8.610 ;
        RECT 24.210 -8.610 25.360 -8.530 ;
        RECT 30.270 -8.230 31.420 -8.150 ;
        RECT 37.710 -8.150 38.160 -8.050 ;
        RECT 44.470 -5.100 44.920 -5.000 ;
        RECT 51.210 -5.000 52.360 -4.920 ;
        RECT 57.270 -4.620 58.420 -4.540 ;
        RECT 64.710 -4.540 65.160 -4.440 ;
        RECT 71.470 -1.490 71.920 -1.390 ;
        RECT 78.210 -1.390 79.360 -1.310 ;
        RECT 84.270 -1.010 85.420 -0.930 ;
        RECT 91.710 -0.930 92.160 -0.830 ;
        RECT 98.470 2.120 98.920 2.220 ;
        RECT 105.210 2.220 106.360 2.300 ;
        RECT 111.270 2.600 112.420 2.680 ;
        RECT 118.710 2.680 119.160 2.780 ;
        RECT 125.470 5.730 125.920 5.830 ;
        RECT 132.210 5.830 133.360 5.910 ;
        RECT 138.270 6.210 139.420 6.290 ;
        RECT 145.710 6.290 146.160 6.390 ;
        RECT 152.470 9.340 152.920 9.440 ;
        RECT 159.210 9.440 160.360 9.520 ;
        RECT 165.270 9.820 166.420 9.900 ;
        RECT 172.710 9.900 173.160 10.000 ;
        RECT 179.470 12.950 179.920 13.050 ;
        RECT 186.210 13.050 187.360 13.130 ;
        RECT 192.270 13.430 193.420 13.510 ;
        RECT 199.710 13.510 200.160 13.610 ;
        RECT 206.470 16.560 206.920 16.660 ;
        RECT 213.210 16.660 214.360 16.740 ;
        RECT 213.210 16.560 213.660 16.660 ;
        RECT 206.470 15.410 206.910 16.560 ;
        RECT 213.220 15.410 213.660 16.560 ;
        RECT 206.470 14.760 207.620 15.410 ;
        RECT 212.510 14.760 213.660 15.410 ;
        RECT 206.470 13.610 206.910 14.760 ;
        RECT 213.220 13.610 213.660 14.760 ;
        RECT 206.470 13.510 206.920 13.610 ;
        RECT 193.670 13.430 194.080 13.490 ;
        RECT 192.270 13.130 194.080 13.430 ;
        RECT 192.270 13.050 193.420 13.130 ;
        RECT 193.670 13.070 194.080 13.130 ;
        RECT 199.050 13.430 199.460 13.490 ;
        RECT 199.710 13.430 200.860 13.510 ;
        RECT 199.050 13.130 200.860 13.430 ;
        RECT 199.050 13.070 199.460 13.130 ;
        RECT 186.210 12.950 186.660 13.050 ;
        RECT 179.470 11.800 179.910 12.950 ;
        RECT 186.220 11.800 186.660 12.950 ;
        RECT 179.470 11.150 180.620 11.800 ;
        RECT 185.510 11.150 186.660 11.800 ;
        RECT 179.470 10.000 179.910 11.150 ;
        RECT 186.220 10.000 186.660 11.150 ;
        RECT 179.470 9.900 179.920 10.000 ;
        RECT 166.670 9.820 167.080 9.880 ;
        RECT 165.270 9.520 167.080 9.820 ;
        RECT 165.270 9.440 166.420 9.520 ;
        RECT 166.670 9.460 167.080 9.520 ;
        RECT 172.050 9.820 172.460 9.880 ;
        RECT 172.710 9.820 173.860 9.900 ;
        RECT 172.050 9.520 173.860 9.820 ;
        RECT 172.050 9.460 172.460 9.520 ;
        RECT 159.210 9.340 159.660 9.440 ;
        RECT 152.470 8.190 152.910 9.340 ;
        RECT 159.220 8.190 159.660 9.340 ;
        RECT 152.470 7.540 153.620 8.190 ;
        RECT 158.510 7.540 159.660 8.190 ;
        RECT 152.470 6.390 152.910 7.540 ;
        RECT 159.220 6.390 159.660 7.540 ;
        RECT 152.470 6.290 152.920 6.390 ;
        RECT 139.670 6.210 140.080 6.270 ;
        RECT 138.270 5.910 140.080 6.210 ;
        RECT 138.270 5.830 139.420 5.910 ;
        RECT 139.670 5.850 140.080 5.910 ;
        RECT 145.050 6.210 145.460 6.270 ;
        RECT 145.710 6.210 146.860 6.290 ;
        RECT 145.050 5.910 146.860 6.210 ;
        RECT 145.050 5.850 145.460 5.910 ;
        RECT 132.210 5.730 132.660 5.830 ;
        RECT 125.470 4.580 125.910 5.730 ;
        RECT 132.220 4.580 132.660 5.730 ;
        RECT 125.470 3.930 126.620 4.580 ;
        RECT 131.510 3.930 132.660 4.580 ;
        RECT 125.470 2.780 125.910 3.930 ;
        RECT 132.220 2.780 132.660 3.930 ;
        RECT 125.470 2.680 125.920 2.780 ;
        RECT 112.670 2.600 113.080 2.660 ;
        RECT 111.270 2.300 113.080 2.600 ;
        RECT 111.270 2.220 112.420 2.300 ;
        RECT 112.670 2.240 113.080 2.300 ;
        RECT 118.050 2.600 118.460 2.660 ;
        RECT 118.710 2.600 119.860 2.680 ;
        RECT 118.050 2.300 119.860 2.600 ;
        RECT 118.050 2.240 118.460 2.300 ;
        RECT 105.210 2.120 105.660 2.220 ;
        RECT 98.470 0.970 98.910 2.120 ;
        RECT 105.220 0.970 105.660 2.120 ;
        RECT 98.470 0.320 99.620 0.970 ;
        RECT 104.510 0.320 105.660 0.970 ;
        RECT 98.470 -0.830 98.910 0.320 ;
        RECT 105.220 -0.830 105.660 0.320 ;
        RECT 98.470 -0.930 98.920 -0.830 ;
        RECT 85.670 -1.010 86.080 -0.950 ;
        RECT 84.270 -1.310 86.080 -1.010 ;
        RECT 84.270 -1.390 85.420 -1.310 ;
        RECT 85.670 -1.370 86.080 -1.310 ;
        RECT 91.050 -1.010 91.460 -0.950 ;
        RECT 91.710 -1.010 92.860 -0.930 ;
        RECT 91.050 -1.310 92.860 -1.010 ;
        RECT 91.050 -1.370 91.460 -1.310 ;
        RECT 78.210 -1.490 78.660 -1.390 ;
        RECT 71.470 -2.640 71.910 -1.490 ;
        RECT 78.220 -2.640 78.660 -1.490 ;
        RECT 71.470 -3.290 72.620 -2.640 ;
        RECT 77.510 -3.290 78.660 -2.640 ;
        RECT 71.470 -4.440 71.910 -3.290 ;
        RECT 78.220 -4.440 78.660 -3.290 ;
        RECT 71.470 -4.540 71.920 -4.440 ;
        RECT 58.670 -4.620 59.080 -4.560 ;
        RECT 57.270 -4.920 59.080 -4.620 ;
        RECT 57.270 -5.000 58.420 -4.920 ;
        RECT 58.670 -4.980 59.080 -4.920 ;
        RECT 64.050 -4.620 64.460 -4.560 ;
        RECT 64.710 -4.620 65.860 -4.540 ;
        RECT 64.050 -4.920 65.860 -4.620 ;
        RECT 64.050 -4.980 64.460 -4.920 ;
        RECT 51.210 -5.100 51.660 -5.000 ;
        RECT 44.470 -6.250 44.910 -5.100 ;
        RECT 51.220 -6.250 51.660 -5.100 ;
        RECT 44.470 -6.900 45.620 -6.250 ;
        RECT 50.510 -6.900 51.660 -6.250 ;
        RECT 44.470 -8.050 44.910 -6.900 ;
        RECT 51.220 -8.050 51.660 -6.900 ;
        RECT 44.470 -8.150 44.920 -8.050 ;
        RECT 31.670 -8.230 32.080 -8.170 ;
        RECT 30.270 -8.530 32.080 -8.230 ;
        RECT 30.270 -8.610 31.420 -8.530 ;
        RECT 31.670 -8.590 32.080 -8.530 ;
        RECT 37.050 -8.230 37.460 -8.170 ;
        RECT 37.710 -8.230 38.860 -8.150 ;
        RECT 37.050 -8.530 38.860 -8.230 ;
        RECT 37.050 -8.590 37.460 -8.530 ;
        RECT 24.210 -8.710 24.660 -8.610 ;
        RECT 17.470 -9.860 17.910 -8.710 ;
        RECT 24.220 -9.860 24.660 -8.710 ;
        RECT 17.470 -10.510 18.620 -9.860 ;
        RECT 23.510 -10.510 24.660 -9.860 ;
        RECT 17.470 -11.660 17.910 -10.510 ;
        RECT 24.220 -11.660 24.660 -10.510 ;
        RECT 17.470 -11.760 17.920 -11.660 ;
        RECT 4.670 -11.840 5.080 -11.780 ;
        RECT 3.270 -12.140 5.080 -11.840 ;
        RECT 3.270 -12.220 4.420 -12.140 ;
        RECT 4.670 -12.200 5.080 -12.140 ;
        RECT 10.050 -11.840 10.460 -11.780 ;
        RECT 10.710 -11.840 11.860 -11.760 ;
        RECT 10.050 -12.140 11.860 -11.840 ;
        RECT 10.050 -12.200 10.460 -12.140 ;
        RECT 3.970 -12.320 4.420 -12.220 ;
        RECT 10.710 -12.220 11.860 -12.140 ;
        RECT 16.770 -11.840 17.920 -11.760 ;
        RECT 24.210 -11.760 24.660 -11.660 ;
        RECT 30.970 -8.710 31.420 -8.610 ;
        RECT 37.710 -8.610 38.860 -8.530 ;
        RECT 43.770 -8.230 44.920 -8.150 ;
        RECT 51.210 -8.150 51.660 -8.050 ;
        RECT 57.970 -5.100 58.420 -5.000 ;
        RECT 64.710 -5.000 65.860 -4.920 ;
        RECT 70.770 -4.620 71.920 -4.540 ;
        RECT 78.210 -4.540 78.660 -4.440 ;
        RECT 84.970 -1.490 85.420 -1.390 ;
        RECT 91.710 -1.390 92.860 -1.310 ;
        RECT 97.770 -1.010 98.920 -0.930 ;
        RECT 105.210 -0.930 105.660 -0.830 ;
        RECT 111.970 2.120 112.420 2.220 ;
        RECT 118.710 2.220 119.860 2.300 ;
        RECT 124.770 2.600 125.920 2.680 ;
        RECT 132.210 2.680 132.660 2.780 ;
        RECT 138.970 5.730 139.420 5.830 ;
        RECT 145.710 5.830 146.860 5.910 ;
        RECT 151.770 6.210 152.920 6.290 ;
        RECT 159.210 6.290 159.660 6.390 ;
        RECT 165.970 9.340 166.420 9.440 ;
        RECT 172.710 9.440 173.860 9.520 ;
        RECT 178.770 9.820 179.920 9.900 ;
        RECT 186.210 9.900 186.660 10.000 ;
        RECT 192.970 12.950 193.420 13.050 ;
        RECT 199.710 13.050 200.860 13.130 ;
        RECT 205.770 13.430 206.920 13.510 ;
        RECT 213.210 13.510 213.660 13.610 ;
        RECT 207.170 13.430 207.580 13.490 ;
        RECT 205.770 13.130 207.580 13.430 ;
        RECT 205.770 13.050 206.920 13.130 ;
        RECT 207.170 13.070 207.580 13.130 ;
        RECT 212.550 13.430 212.960 13.490 ;
        RECT 213.210 13.430 214.360 13.510 ;
        RECT 212.550 13.130 214.360 13.430 ;
        RECT 212.550 13.070 212.960 13.130 ;
        RECT 199.710 12.950 200.160 13.050 ;
        RECT 192.970 11.800 193.410 12.950 ;
        RECT 199.720 11.800 200.160 12.950 ;
        RECT 192.970 11.150 194.120 11.800 ;
        RECT 199.010 11.150 200.160 11.800 ;
        RECT 192.970 10.000 193.410 11.150 ;
        RECT 199.720 10.000 200.160 11.150 ;
        RECT 192.970 9.900 193.420 10.000 ;
        RECT 180.170 9.820 180.580 9.880 ;
        RECT 178.770 9.520 180.580 9.820 ;
        RECT 178.770 9.440 179.920 9.520 ;
        RECT 180.170 9.460 180.580 9.520 ;
        RECT 185.550 9.820 185.960 9.880 ;
        RECT 186.210 9.820 187.360 9.900 ;
        RECT 185.550 9.520 187.360 9.820 ;
        RECT 185.550 9.460 185.960 9.520 ;
        RECT 172.710 9.340 173.160 9.440 ;
        RECT 165.970 8.190 166.410 9.340 ;
        RECT 172.720 8.190 173.160 9.340 ;
        RECT 165.970 7.540 167.120 8.190 ;
        RECT 172.010 7.540 173.160 8.190 ;
        RECT 165.970 6.390 166.410 7.540 ;
        RECT 172.720 6.390 173.160 7.540 ;
        RECT 165.970 6.290 166.420 6.390 ;
        RECT 153.170 6.210 153.580 6.270 ;
        RECT 151.770 5.910 153.580 6.210 ;
        RECT 151.770 5.830 152.920 5.910 ;
        RECT 153.170 5.850 153.580 5.910 ;
        RECT 158.550 6.210 158.960 6.270 ;
        RECT 159.210 6.210 160.360 6.290 ;
        RECT 158.550 5.910 160.360 6.210 ;
        RECT 158.550 5.850 158.960 5.910 ;
        RECT 145.710 5.730 146.160 5.830 ;
        RECT 138.970 4.580 139.410 5.730 ;
        RECT 145.720 4.580 146.160 5.730 ;
        RECT 138.970 3.930 140.120 4.580 ;
        RECT 145.010 3.930 146.160 4.580 ;
        RECT 138.970 2.780 139.410 3.930 ;
        RECT 145.720 2.780 146.160 3.930 ;
        RECT 138.970 2.680 139.420 2.780 ;
        RECT 126.170 2.600 126.580 2.660 ;
        RECT 124.770 2.300 126.580 2.600 ;
        RECT 124.770 2.220 125.920 2.300 ;
        RECT 126.170 2.240 126.580 2.300 ;
        RECT 131.550 2.600 131.960 2.660 ;
        RECT 132.210 2.600 133.360 2.680 ;
        RECT 131.550 2.300 133.360 2.600 ;
        RECT 131.550 2.240 131.960 2.300 ;
        RECT 118.710 2.120 119.160 2.220 ;
        RECT 111.970 0.970 112.410 2.120 ;
        RECT 118.720 0.970 119.160 2.120 ;
        RECT 111.970 0.320 113.120 0.970 ;
        RECT 118.010 0.320 119.160 0.970 ;
        RECT 111.970 -0.830 112.410 0.320 ;
        RECT 118.720 -0.830 119.160 0.320 ;
        RECT 111.970 -0.930 112.420 -0.830 ;
        RECT 99.170 -1.010 99.580 -0.950 ;
        RECT 97.770 -1.310 99.580 -1.010 ;
        RECT 97.770 -1.390 98.920 -1.310 ;
        RECT 99.170 -1.370 99.580 -1.310 ;
        RECT 104.550 -1.010 104.960 -0.950 ;
        RECT 105.210 -1.010 106.360 -0.930 ;
        RECT 104.550 -1.310 106.360 -1.010 ;
        RECT 104.550 -1.370 104.960 -1.310 ;
        RECT 91.710 -1.490 92.160 -1.390 ;
        RECT 84.970 -2.640 85.410 -1.490 ;
        RECT 91.720 -2.640 92.160 -1.490 ;
        RECT 84.970 -3.290 86.120 -2.640 ;
        RECT 91.010 -3.290 92.160 -2.640 ;
        RECT 84.970 -4.440 85.410 -3.290 ;
        RECT 91.720 -4.440 92.160 -3.290 ;
        RECT 84.970 -4.540 85.420 -4.440 ;
        RECT 72.170 -4.620 72.580 -4.560 ;
        RECT 70.770 -4.920 72.580 -4.620 ;
        RECT 70.770 -5.000 71.920 -4.920 ;
        RECT 72.170 -4.980 72.580 -4.920 ;
        RECT 77.550 -4.620 77.960 -4.560 ;
        RECT 78.210 -4.620 79.360 -4.540 ;
        RECT 77.550 -4.920 79.360 -4.620 ;
        RECT 77.550 -4.980 77.960 -4.920 ;
        RECT 64.710 -5.100 65.160 -5.000 ;
        RECT 57.970 -6.250 58.410 -5.100 ;
        RECT 64.720 -6.250 65.160 -5.100 ;
        RECT 57.970 -6.900 59.120 -6.250 ;
        RECT 64.010 -6.900 65.160 -6.250 ;
        RECT 57.970 -8.050 58.410 -6.900 ;
        RECT 64.720 -8.050 65.160 -6.900 ;
        RECT 57.970 -8.150 58.420 -8.050 ;
        RECT 45.170 -8.230 45.580 -8.170 ;
        RECT 43.770 -8.530 45.580 -8.230 ;
        RECT 43.770 -8.610 44.920 -8.530 ;
        RECT 45.170 -8.590 45.580 -8.530 ;
        RECT 50.550 -8.230 50.960 -8.170 ;
        RECT 51.210 -8.230 52.360 -8.150 ;
        RECT 50.550 -8.530 52.360 -8.230 ;
        RECT 50.550 -8.590 50.960 -8.530 ;
        RECT 37.710 -8.710 38.160 -8.610 ;
        RECT 30.970 -9.860 31.410 -8.710 ;
        RECT 37.720 -9.860 38.160 -8.710 ;
        RECT 30.970 -10.510 32.120 -9.860 ;
        RECT 37.010 -10.510 38.160 -9.860 ;
        RECT 30.970 -11.660 31.410 -10.510 ;
        RECT 37.720 -11.660 38.160 -10.510 ;
        RECT 30.970 -11.760 31.420 -11.660 ;
        RECT 18.170 -11.840 18.580 -11.780 ;
        RECT 16.770 -12.140 18.580 -11.840 ;
        RECT 16.770 -12.220 17.920 -12.140 ;
        RECT 18.170 -12.200 18.580 -12.140 ;
        RECT 23.550 -11.840 23.960 -11.780 ;
        RECT 24.210 -11.840 25.360 -11.760 ;
        RECT 23.550 -12.140 25.360 -11.840 ;
        RECT 23.550 -12.200 23.960 -12.140 ;
        RECT 10.710 -12.320 11.160 -12.220 ;
        RECT 3.970 -13.470 4.410 -12.320 ;
        RECT 10.720 -13.470 11.160 -12.320 ;
        RECT 3.970 -14.120 5.120 -13.470 ;
        RECT 10.010 -14.120 11.160 -13.470 ;
        RECT 3.970 -15.270 4.410 -14.120 ;
        RECT 10.720 -15.270 11.160 -14.120 ;
        RECT 3.970 -15.370 4.420 -15.270 ;
        RECT 3.270 -15.450 4.420 -15.370 ;
        RECT 10.710 -15.370 11.160 -15.270 ;
        RECT 17.470 -12.320 17.920 -12.220 ;
        RECT 24.210 -12.220 25.360 -12.140 ;
        RECT 30.270 -11.840 31.420 -11.760 ;
        RECT 37.710 -11.760 38.160 -11.660 ;
        RECT 44.470 -8.710 44.920 -8.610 ;
        RECT 51.210 -8.610 52.360 -8.530 ;
        RECT 57.270 -8.230 58.420 -8.150 ;
        RECT 64.710 -8.150 65.160 -8.050 ;
        RECT 71.470 -5.100 71.920 -5.000 ;
        RECT 78.210 -5.000 79.360 -4.920 ;
        RECT 84.270 -4.620 85.420 -4.540 ;
        RECT 91.710 -4.540 92.160 -4.440 ;
        RECT 98.470 -1.490 98.920 -1.390 ;
        RECT 105.210 -1.390 106.360 -1.310 ;
        RECT 111.270 -1.010 112.420 -0.930 ;
        RECT 118.710 -0.930 119.160 -0.830 ;
        RECT 125.470 2.120 125.920 2.220 ;
        RECT 132.210 2.220 133.360 2.300 ;
        RECT 138.270 2.600 139.420 2.680 ;
        RECT 145.710 2.680 146.160 2.780 ;
        RECT 152.470 5.730 152.920 5.830 ;
        RECT 159.210 5.830 160.360 5.910 ;
        RECT 165.270 6.210 166.420 6.290 ;
        RECT 172.710 6.290 173.160 6.390 ;
        RECT 179.470 9.340 179.920 9.440 ;
        RECT 186.210 9.440 187.360 9.520 ;
        RECT 192.270 9.820 193.420 9.900 ;
        RECT 199.710 9.900 200.160 10.000 ;
        RECT 206.470 12.950 206.920 13.050 ;
        RECT 213.210 13.050 214.360 13.130 ;
        RECT 213.210 12.950 213.660 13.050 ;
        RECT 206.470 11.800 206.910 12.950 ;
        RECT 213.220 11.800 213.660 12.950 ;
        RECT 206.470 11.150 207.620 11.800 ;
        RECT 212.510 11.150 213.660 11.800 ;
        RECT 206.470 10.000 206.910 11.150 ;
        RECT 213.220 10.000 213.660 11.150 ;
        RECT 206.470 9.900 206.920 10.000 ;
        RECT 193.670 9.820 194.080 9.880 ;
        RECT 192.270 9.520 194.080 9.820 ;
        RECT 192.270 9.440 193.420 9.520 ;
        RECT 193.670 9.460 194.080 9.520 ;
        RECT 199.050 9.820 199.460 9.880 ;
        RECT 199.710 9.820 200.860 9.900 ;
        RECT 199.050 9.520 200.860 9.820 ;
        RECT 199.050 9.460 199.460 9.520 ;
        RECT 186.210 9.340 186.660 9.440 ;
        RECT 179.470 8.190 179.910 9.340 ;
        RECT 186.220 8.190 186.660 9.340 ;
        RECT 179.470 7.540 180.620 8.190 ;
        RECT 185.510 7.540 186.660 8.190 ;
        RECT 179.470 6.390 179.910 7.540 ;
        RECT 186.220 6.390 186.660 7.540 ;
        RECT 179.470 6.290 179.920 6.390 ;
        RECT 166.670 6.210 167.080 6.270 ;
        RECT 165.270 5.910 167.080 6.210 ;
        RECT 165.270 5.830 166.420 5.910 ;
        RECT 166.670 5.850 167.080 5.910 ;
        RECT 172.050 6.210 172.460 6.270 ;
        RECT 172.710 6.210 173.860 6.290 ;
        RECT 172.050 5.910 173.860 6.210 ;
        RECT 172.050 5.850 172.460 5.910 ;
        RECT 159.210 5.730 159.660 5.830 ;
        RECT 152.470 4.580 152.910 5.730 ;
        RECT 159.220 4.580 159.660 5.730 ;
        RECT 152.470 3.930 153.620 4.580 ;
        RECT 158.510 3.930 159.660 4.580 ;
        RECT 152.470 2.780 152.910 3.930 ;
        RECT 159.220 2.780 159.660 3.930 ;
        RECT 152.470 2.680 152.920 2.780 ;
        RECT 139.670 2.600 140.080 2.660 ;
        RECT 138.270 2.300 140.080 2.600 ;
        RECT 138.270 2.220 139.420 2.300 ;
        RECT 139.670 2.240 140.080 2.300 ;
        RECT 145.050 2.600 145.460 2.660 ;
        RECT 145.710 2.600 146.860 2.680 ;
        RECT 145.050 2.300 146.860 2.600 ;
        RECT 145.050 2.240 145.460 2.300 ;
        RECT 132.210 2.120 132.660 2.220 ;
        RECT 125.470 0.970 125.910 2.120 ;
        RECT 132.220 0.970 132.660 2.120 ;
        RECT 125.470 0.320 126.620 0.970 ;
        RECT 131.510 0.320 132.660 0.970 ;
        RECT 125.470 -0.830 125.910 0.320 ;
        RECT 132.220 -0.830 132.660 0.320 ;
        RECT 125.470 -0.930 125.920 -0.830 ;
        RECT 112.670 -1.010 113.080 -0.950 ;
        RECT 111.270 -1.310 113.080 -1.010 ;
        RECT 111.270 -1.390 112.420 -1.310 ;
        RECT 112.670 -1.370 113.080 -1.310 ;
        RECT 118.050 -1.010 118.460 -0.950 ;
        RECT 118.710 -1.010 119.860 -0.930 ;
        RECT 118.050 -1.310 119.860 -1.010 ;
        RECT 118.050 -1.370 118.460 -1.310 ;
        RECT 105.210 -1.490 105.660 -1.390 ;
        RECT 98.470 -2.640 98.910 -1.490 ;
        RECT 105.220 -2.640 105.660 -1.490 ;
        RECT 98.470 -3.290 99.620 -2.640 ;
        RECT 104.510 -3.290 105.660 -2.640 ;
        RECT 98.470 -4.440 98.910 -3.290 ;
        RECT 105.220 -4.440 105.660 -3.290 ;
        RECT 98.470 -4.540 98.920 -4.440 ;
        RECT 85.670 -4.620 86.080 -4.560 ;
        RECT 84.270 -4.920 86.080 -4.620 ;
        RECT 84.270 -5.000 85.420 -4.920 ;
        RECT 85.670 -4.980 86.080 -4.920 ;
        RECT 91.050 -4.620 91.460 -4.560 ;
        RECT 91.710 -4.620 92.860 -4.540 ;
        RECT 91.050 -4.920 92.860 -4.620 ;
        RECT 91.050 -4.980 91.460 -4.920 ;
        RECT 78.210 -5.100 78.660 -5.000 ;
        RECT 71.470 -6.250 71.910 -5.100 ;
        RECT 78.220 -6.250 78.660 -5.100 ;
        RECT 71.470 -6.900 72.620 -6.250 ;
        RECT 77.510 -6.900 78.660 -6.250 ;
        RECT 71.470 -8.050 71.910 -6.900 ;
        RECT 78.220 -8.050 78.660 -6.900 ;
        RECT 71.470 -8.150 71.920 -8.050 ;
        RECT 58.670 -8.230 59.080 -8.170 ;
        RECT 57.270 -8.530 59.080 -8.230 ;
        RECT 57.270 -8.610 58.420 -8.530 ;
        RECT 58.670 -8.590 59.080 -8.530 ;
        RECT 64.050 -8.230 64.460 -8.170 ;
        RECT 64.710 -8.230 65.860 -8.150 ;
        RECT 64.050 -8.530 65.860 -8.230 ;
        RECT 64.050 -8.590 64.460 -8.530 ;
        RECT 51.210 -8.710 51.660 -8.610 ;
        RECT 44.470 -9.860 44.910 -8.710 ;
        RECT 51.220 -9.860 51.660 -8.710 ;
        RECT 44.470 -10.510 45.620 -9.860 ;
        RECT 50.510 -10.510 51.660 -9.860 ;
        RECT 44.470 -11.660 44.910 -10.510 ;
        RECT 51.220 -11.660 51.660 -10.510 ;
        RECT 44.470 -11.760 44.920 -11.660 ;
        RECT 31.670 -11.840 32.080 -11.780 ;
        RECT 30.270 -12.140 32.080 -11.840 ;
        RECT 30.270 -12.220 31.420 -12.140 ;
        RECT 31.670 -12.200 32.080 -12.140 ;
        RECT 37.050 -11.840 37.460 -11.780 ;
        RECT 37.710 -11.840 38.860 -11.760 ;
        RECT 37.050 -12.140 38.860 -11.840 ;
        RECT 37.050 -12.200 37.460 -12.140 ;
        RECT 24.210 -12.320 24.660 -12.220 ;
        RECT 17.470 -13.470 17.910 -12.320 ;
        RECT 24.220 -13.470 24.660 -12.320 ;
        RECT 17.470 -14.120 18.620 -13.470 ;
        RECT 23.510 -14.120 24.660 -13.470 ;
        RECT 17.470 -15.270 17.910 -14.120 ;
        RECT 24.220 -15.270 24.660 -14.120 ;
        RECT 17.470 -15.370 17.920 -15.270 ;
        RECT 4.670 -15.450 5.080 -15.390 ;
        RECT 3.270 -15.750 5.080 -15.450 ;
        RECT 3.270 -15.830 4.420 -15.750 ;
        RECT 4.670 -15.810 5.080 -15.750 ;
        RECT 10.050 -15.450 10.460 -15.390 ;
        RECT 10.710 -15.450 11.860 -15.370 ;
        RECT 10.050 -15.750 11.860 -15.450 ;
        RECT 10.050 -15.810 10.460 -15.750 ;
        RECT 3.970 -15.930 4.420 -15.830 ;
        RECT 10.710 -15.830 11.860 -15.750 ;
        RECT 16.770 -15.450 17.920 -15.370 ;
        RECT 24.210 -15.370 24.660 -15.270 ;
        RECT 30.970 -12.320 31.420 -12.220 ;
        RECT 37.710 -12.220 38.860 -12.140 ;
        RECT 43.770 -11.840 44.920 -11.760 ;
        RECT 51.210 -11.760 51.660 -11.660 ;
        RECT 57.970 -8.710 58.420 -8.610 ;
        RECT 64.710 -8.610 65.860 -8.530 ;
        RECT 70.770 -8.230 71.920 -8.150 ;
        RECT 78.210 -8.150 78.660 -8.050 ;
        RECT 84.970 -5.100 85.420 -5.000 ;
        RECT 91.710 -5.000 92.860 -4.920 ;
        RECT 97.770 -4.620 98.920 -4.540 ;
        RECT 105.210 -4.540 105.660 -4.440 ;
        RECT 111.970 -1.490 112.420 -1.390 ;
        RECT 118.710 -1.390 119.860 -1.310 ;
        RECT 124.770 -1.010 125.920 -0.930 ;
        RECT 132.210 -0.930 132.660 -0.830 ;
        RECT 138.970 2.120 139.420 2.220 ;
        RECT 145.710 2.220 146.860 2.300 ;
        RECT 151.770 2.600 152.920 2.680 ;
        RECT 159.210 2.680 159.660 2.780 ;
        RECT 165.970 5.730 166.420 5.830 ;
        RECT 172.710 5.830 173.860 5.910 ;
        RECT 178.770 6.210 179.920 6.290 ;
        RECT 186.210 6.290 186.660 6.390 ;
        RECT 192.970 9.340 193.420 9.440 ;
        RECT 199.710 9.440 200.860 9.520 ;
        RECT 205.770 9.820 206.920 9.900 ;
        RECT 213.210 9.900 213.660 10.000 ;
        RECT 207.170 9.820 207.580 9.880 ;
        RECT 205.770 9.520 207.580 9.820 ;
        RECT 205.770 9.440 206.920 9.520 ;
        RECT 207.170 9.460 207.580 9.520 ;
        RECT 212.550 9.820 212.960 9.880 ;
        RECT 213.210 9.820 214.360 9.900 ;
        RECT 212.550 9.520 214.360 9.820 ;
        RECT 212.550 9.460 212.960 9.520 ;
        RECT 199.710 9.340 200.160 9.440 ;
        RECT 192.970 8.190 193.410 9.340 ;
        RECT 199.720 8.190 200.160 9.340 ;
        RECT 192.970 7.540 194.120 8.190 ;
        RECT 199.010 7.540 200.160 8.190 ;
        RECT 192.970 6.390 193.410 7.540 ;
        RECT 199.720 6.390 200.160 7.540 ;
        RECT 192.970 6.290 193.420 6.390 ;
        RECT 180.170 6.210 180.580 6.270 ;
        RECT 178.770 5.910 180.580 6.210 ;
        RECT 178.770 5.830 179.920 5.910 ;
        RECT 180.170 5.850 180.580 5.910 ;
        RECT 185.550 6.210 185.960 6.270 ;
        RECT 186.210 6.210 187.360 6.290 ;
        RECT 185.550 5.910 187.360 6.210 ;
        RECT 185.550 5.850 185.960 5.910 ;
        RECT 172.710 5.730 173.160 5.830 ;
        RECT 165.970 4.580 166.410 5.730 ;
        RECT 172.720 4.580 173.160 5.730 ;
        RECT 165.970 3.930 167.120 4.580 ;
        RECT 172.010 3.930 173.160 4.580 ;
        RECT 165.970 2.780 166.410 3.930 ;
        RECT 172.720 2.780 173.160 3.930 ;
        RECT 165.970 2.680 166.420 2.780 ;
        RECT 153.170 2.600 153.580 2.660 ;
        RECT 151.770 2.300 153.580 2.600 ;
        RECT 151.770 2.220 152.920 2.300 ;
        RECT 153.170 2.240 153.580 2.300 ;
        RECT 158.550 2.600 158.960 2.660 ;
        RECT 159.210 2.600 160.360 2.680 ;
        RECT 158.550 2.300 160.360 2.600 ;
        RECT 158.550 2.240 158.960 2.300 ;
        RECT 145.710 2.120 146.160 2.220 ;
        RECT 138.970 0.970 139.410 2.120 ;
        RECT 145.720 0.970 146.160 2.120 ;
        RECT 138.970 0.320 140.120 0.970 ;
        RECT 145.010 0.320 146.160 0.970 ;
        RECT 138.970 -0.830 139.410 0.320 ;
        RECT 145.720 -0.830 146.160 0.320 ;
        RECT 138.970 -0.930 139.420 -0.830 ;
        RECT 126.170 -1.010 126.580 -0.950 ;
        RECT 124.770 -1.310 126.580 -1.010 ;
        RECT 124.770 -1.390 125.920 -1.310 ;
        RECT 126.170 -1.370 126.580 -1.310 ;
        RECT 131.550 -1.010 131.960 -0.950 ;
        RECT 132.210 -1.010 133.360 -0.930 ;
        RECT 131.550 -1.310 133.360 -1.010 ;
        RECT 131.550 -1.370 131.960 -1.310 ;
        RECT 118.710 -1.490 119.160 -1.390 ;
        RECT 111.970 -2.640 112.410 -1.490 ;
        RECT 118.720 -2.640 119.160 -1.490 ;
        RECT 111.970 -3.290 113.120 -2.640 ;
        RECT 118.010 -3.290 119.160 -2.640 ;
        RECT 111.970 -4.440 112.410 -3.290 ;
        RECT 118.720 -4.440 119.160 -3.290 ;
        RECT 111.970 -4.540 112.420 -4.440 ;
        RECT 99.170 -4.620 99.580 -4.560 ;
        RECT 97.770 -4.920 99.580 -4.620 ;
        RECT 97.770 -5.000 98.920 -4.920 ;
        RECT 99.170 -4.980 99.580 -4.920 ;
        RECT 104.550 -4.620 104.960 -4.560 ;
        RECT 105.210 -4.620 106.360 -4.540 ;
        RECT 104.550 -4.920 106.360 -4.620 ;
        RECT 104.550 -4.980 104.960 -4.920 ;
        RECT 91.710 -5.100 92.160 -5.000 ;
        RECT 84.970 -6.250 85.410 -5.100 ;
        RECT 91.720 -6.250 92.160 -5.100 ;
        RECT 84.970 -6.900 86.120 -6.250 ;
        RECT 91.010 -6.900 92.160 -6.250 ;
        RECT 84.970 -8.050 85.410 -6.900 ;
        RECT 91.720 -8.050 92.160 -6.900 ;
        RECT 84.970 -8.150 85.420 -8.050 ;
        RECT 72.170 -8.230 72.580 -8.170 ;
        RECT 70.770 -8.530 72.580 -8.230 ;
        RECT 70.770 -8.610 71.920 -8.530 ;
        RECT 72.170 -8.590 72.580 -8.530 ;
        RECT 77.550 -8.230 77.960 -8.170 ;
        RECT 78.210 -8.230 79.360 -8.150 ;
        RECT 77.550 -8.530 79.360 -8.230 ;
        RECT 77.550 -8.590 77.960 -8.530 ;
        RECT 64.710 -8.710 65.160 -8.610 ;
        RECT 57.970 -9.860 58.410 -8.710 ;
        RECT 64.720 -9.860 65.160 -8.710 ;
        RECT 57.970 -10.510 59.120 -9.860 ;
        RECT 64.010 -10.510 65.160 -9.860 ;
        RECT 57.970 -11.660 58.410 -10.510 ;
        RECT 64.720 -11.660 65.160 -10.510 ;
        RECT 57.970 -11.760 58.420 -11.660 ;
        RECT 45.170 -11.840 45.580 -11.780 ;
        RECT 43.770 -12.140 45.580 -11.840 ;
        RECT 43.770 -12.220 44.920 -12.140 ;
        RECT 45.170 -12.200 45.580 -12.140 ;
        RECT 50.550 -11.840 50.960 -11.780 ;
        RECT 51.210 -11.840 52.360 -11.760 ;
        RECT 50.550 -12.140 52.360 -11.840 ;
        RECT 50.550 -12.200 50.960 -12.140 ;
        RECT 37.710 -12.320 38.160 -12.220 ;
        RECT 30.970 -13.470 31.410 -12.320 ;
        RECT 37.720 -13.470 38.160 -12.320 ;
        RECT 30.970 -14.120 32.120 -13.470 ;
        RECT 37.010 -14.120 38.160 -13.470 ;
        RECT 30.970 -15.270 31.410 -14.120 ;
        RECT 37.720 -15.270 38.160 -14.120 ;
        RECT 30.970 -15.370 31.420 -15.270 ;
        RECT 18.170 -15.450 18.580 -15.390 ;
        RECT 16.770 -15.750 18.580 -15.450 ;
        RECT 16.770 -15.830 17.920 -15.750 ;
        RECT 18.170 -15.810 18.580 -15.750 ;
        RECT 23.550 -15.450 23.960 -15.390 ;
        RECT 24.210 -15.450 25.360 -15.370 ;
        RECT 23.550 -15.750 25.360 -15.450 ;
        RECT 23.550 -15.810 23.960 -15.750 ;
        RECT 10.710 -15.930 11.160 -15.830 ;
        RECT 3.970 -17.080 4.410 -15.930 ;
        RECT 10.720 -17.080 11.160 -15.930 ;
        RECT 3.970 -17.730 5.120 -17.080 ;
        RECT 10.010 -17.730 11.160 -17.080 ;
        RECT 3.970 -18.880 4.410 -17.730 ;
        RECT 10.720 -18.880 11.160 -17.730 ;
        RECT 3.970 -18.980 4.420 -18.880 ;
        RECT 3.270 -19.060 4.420 -18.980 ;
        RECT 10.710 -18.980 11.160 -18.880 ;
        RECT 17.470 -15.930 17.920 -15.830 ;
        RECT 24.210 -15.830 25.360 -15.750 ;
        RECT 30.270 -15.450 31.420 -15.370 ;
        RECT 37.710 -15.370 38.160 -15.270 ;
        RECT 44.470 -12.320 44.920 -12.220 ;
        RECT 51.210 -12.220 52.360 -12.140 ;
        RECT 57.270 -11.840 58.420 -11.760 ;
        RECT 64.710 -11.760 65.160 -11.660 ;
        RECT 71.470 -8.710 71.920 -8.610 ;
        RECT 78.210 -8.610 79.360 -8.530 ;
        RECT 84.270 -8.230 85.420 -8.150 ;
        RECT 91.710 -8.150 92.160 -8.050 ;
        RECT 98.470 -5.100 98.920 -5.000 ;
        RECT 105.210 -5.000 106.360 -4.920 ;
        RECT 111.270 -4.620 112.420 -4.540 ;
        RECT 118.710 -4.540 119.160 -4.440 ;
        RECT 125.470 -1.490 125.920 -1.390 ;
        RECT 132.210 -1.390 133.360 -1.310 ;
        RECT 138.270 -1.010 139.420 -0.930 ;
        RECT 145.710 -0.930 146.160 -0.830 ;
        RECT 152.470 2.120 152.920 2.220 ;
        RECT 159.210 2.220 160.360 2.300 ;
        RECT 165.270 2.600 166.420 2.680 ;
        RECT 172.710 2.680 173.160 2.780 ;
        RECT 179.470 5.730 179.920 5.830 ;
        RECT 186.210 5.830 187.360 5.910 ;
        RECT 192.270 6.210 193.420 6.290 ;
        RECT 199.710 6.290 200.160 6.390 ;
        RECT 206.470 9.340 206.920 9.440 ;
        RECT 213.210 9.440 214.360 9.520 ;
        RECT 213.210 9.340 213.660 9.440 ;
        RECT 206.470 8.190 206.910 9.340 ;
        RECT 213.220 8.190 213.660 9.340 ;
        RECT 206.470 7.540 207.620 8.190 ;
        RECT 212.510 7.540 213.660 8.190 ;
        RECT 206.470 6.390 206.910 7.540 ;
        RECT 213.220 6.390 213.660 7.540 ;
        RECT 206.470 6.290 206.920 6.390 ;
        RECT 193.670 6.210 194.080 6.270 ;
        RECT 192.270 5.910 194.080 6.210 ;
        RECT 192.270 5.830 193.420 5.910 ;
        RECT 193.670 5.850 194.080 5.910 ;
        RECT 199.050 6.210 199.460 6.270 ;
        RECT 199.710 6.210 200.860 6.290 ;
        RECT 199.050 5.910 200.860 6.210 ;
        RECT 199.050 5.850 199.460 5.910 ;
        RECT 186.210 5.730 186.660 5.830 ;
        RECT 179.470 4.580 179.910 5.730 ;
        RECT 186.220 4.580 186.660 5.730 ;
        RECT 179.470 3.930 180.620 4.580 ;
        RECT 185.510 3.930 186.660 4.580 ;
        RECT 179.470 2.780 179.910 3.930 ;
        RECT 186.220 2.780 186.660 3.930 ;
        RECT 179.470 2.680 179.920 2.780 ;
        RECT 166.670 2.600 167.080 2.660 ;
        RECT 165.270 2.300 167.080 2.600 ;
        RECT 165.270 2.220 166.420 2.300 ;
        RECT 166.670 2.240 167.080 2.300 ;
        RECT 172.050 2.600 172.460 2.660 ;
        RECT 172.710 2.600 173.860 2.680 ;
        RECT 172.050 2.300 173.860 2.600 ;
        RECT 172.050 2.240 172.460 2.300 ;
        RECT 159.210 2.120 159.660 2.220 ;
        RECT 152.470 0.970 152.910 2.120 ;
        RECT 159.220 0.970 159.660 2.120 ;
        RECT 152.470 0.320 153.620 0.970 ;
        RECT 158.510 0.320 159.660 0.970 ;
        RECT 152.470 -0.830 152.910 0.320 ;
        RECT 159.220 -0.830 159.660 0.320 ;
        RECT 152.470 -0.930 152.920 -0.830 ;
        RECT 139.670 -1.010 140.080 -0.950 ;
        RECT 138.270 -1.310 140.080 -1.010 ;
        RECT 138.270 -1.390 139.420 -1.310 ;
        RECT 139.670 -1.370 140.080 -1.310 ;
        RECT 145.050 -1.010 145.460 -0.950 ;
        RECT 145.710 -1.010 146.860 -0.930 ;
        RECT 145.050 -1.310 146.860 -1.010 ;
        RECT 145.050 -1.370 145.460 -1.310 ;
        RECT 132.210 -1.490 132.660 -1.390 ;
        RECT 125.470 -2.640 125.910 -1.490 ;
        RECT 132.220 -2.640 132.660 -1.490 ;
        RECT 125.470 -3.290 126.620 -2.640 ;
        RECT 131.510 -3.290 132.660 -2.640 ;
        RECT 125.470 -4.440 125.910 -3.290 ;
        RECT 132.220 -4.440 132.660 -3.290 ;
        RECT 125.470 -4.540 125.920 -4.440 ;
        RECT 112.670 -4.620 113.080 -4.560 ;
        RECT 111.270 -4.920 113.080 -4.620 ;
        RECT 111.270 -5.000 112.420 -4.920 ;
        RECT 112.670 -4.980 113.080 -4.920 ;
        RECT 118.050 -4.620 118.460 -4.560 ;
        RECT 118.710 -4.620 119.860 -4.540 ;
        RECT 118.050 -4.920 119.860 -4.620 ;
        RECT 118.050 -4.980 118.460 -4.920 ;
        RECT 105.210 -5.100 105.660 -5.000 ;
        RECT 98.470 -6.250 98.910 -5.100 ;
        RECT 105.220 -6.250 105.660 -5.100 ;
        RECT 98.470 -6.900 99.620 -6.250 ;
        RECT 104.510 -6.900 105.660 -6.250 ;
        RECT 98.470 -8.050 98.910 -6.900 ;
        RECT 105.220 -8.050 105.660 -6.900 ;
        RECT 98.470 -8.150 98.920 -8.050 ;
        RECT 85.670 -8.230 86.080 -8.170 ;
        RECT 84.270 -8.530 86.080 -8.230 ;
        RECT 84.270 -8.610 85.420 -8.530 ;
        RECT 85.670 -8.590 86.080 -8.530 ;
        RECT 91.050 -8.230 91.460 -8.170 ;
        RECT 91.710 -8.230 92.860 -8.150 ;
        RECT 91.050 -8.530 92.860 -8.230 ;
        RECT 91.050 -8.590 91.460 -8.530 ;
        RECT 78.210 -8.710 78.660 -8.610 ;
        RECT 71.470 -9.860 71.910 -8.710 ;
        RECT 78.220 -9.860 78.660 -8.710 ;
        RECT 71.470 -10.510 72.620 -9.860 ;
        RECT 77.510 -10.510 78.660 -9.860 ;
        RECT 71.470 -11.660 71.910 -10.510 ;
        RECT 78.220 -11.660 78.660 -10.510 ;
        RECT 71.470 -11.760 71.920 -11.660 ;
        RECT 58.670 -11.840 59.080 -11.780 ;
        RECT 57.270 -12.140 59.080 -11.840 ;
        RECT 57.270 -12.220 58.420 -12.140 ;
        RECT 58.670 -12.200 59.080 -12.140 ;
        RECT 64.050 -11.840 64.460 -11.780 ;
        RECT 64.710 -11.840 65.860 -11.760 ;
        RECT 64.050 -12.140 65.860 -11.840 ;
        RECT 64.050 -12.200 64.460 -12.140 ;
        RECT 51.210 -12.320 51.660 -12.220 ;
        RECT 44.470 -13.470 44.910 -12.320 ;
        RECT 51.220 -13.470 51.660 -12.320 ;
        RECT 44.470 -14.120 45.620 -13.470 ;
        RECT 50.510 -14.120 51.660 -13.470 ;
        RECT 44.470 -15.270 44.910 -14.120 ;
        RECT 51.220 -15.270 51.660 -14.120 ;
        RECT 44.470 -15.370 44.920 -15.270 ;
        RECT 31.670 -15.450 32.080 -15.390 ;
        RECT 30.270 -15.750 32.080 -15.450 ;
        RECT 30.270 -15.830 31.420 -15.750 ;
        RECT 31.670 -15.810 32.080 -15.750 ;
        RECT 37.050 -15.450 37.460 -15.390 ;
        RECT 37.710 -15.450 38.860 -15.370 ;
        RECT 37.050 -15.750 38.860 -15.450 ;
        RECT 37.050 -15.810 37.460 -15.750 ;
        RECT 24.210 -15.930 24.660 -15.830 ;
        RECT 17.470 -17.080 17.910 -15.930 ;
        RECT 24.220 -17.080 24.660 -15.930 ;
        RECT 17.470 -17.730 18.620 -17.080 ;
        RECT 23.510 -17.730 24.660 -17.080 ;
        RECT 17.470 -18.880 17.910 -17.730 ;
        RECT 24.220 -18.880 24.660 -17.730 ;
        RECT 17.470 -18.980 17.920 -18.880 ;
        RECT 4.670 -19.060 5.080 -19.000 ;
        RECT 3.270 -19.360 5.080 -19.060 ;
        RECT 3.270 -19.440 4.420 -19.360 ;
        RECT 4.670 -19.420 5.080 -19.360 ;
        RECT 10.050 -19.060 10.460 -19.000 ;
        RECT 10.710 -19.060 11.860 -18.980 ;
        RECT 10.050 -19.360 11.860 -19.060 ;
        RECT 10.050 -19.420 10.460 -19.360 ;
        RECT 3.970 -19.540 4.420 -19.440 ;
        RECT 10.710 -19.440 11.860 -19.360 ;
        RECT 16.770 -19.060 17.920 -18.980 ;
        RECT 24.210 -18.980 24.660 -18.880 ;
        RECT 30.970 -15.930 31.420 -15.830 ;
        RECT 37.710 -15.830 38.860 -15.750 ;
        RECT 43.770 -15.450 44.920 -15.370 ;
        RECT 51.210 -15.370 51.660 -15.270 ;
        RECT 57.970 -12.320 58.420 -12.220 ;
        RECT 64.710 -12.220 65.860 -12.140 ;
        RECT 70.770 -11.840 71.920 -11.760 ;
        RECT 78.210 -11.760 78.660 -11.660 ;
        RECT 84.970 -8.710 85.420 -8.610 ;
        RECT 91.710 -8.610 92.860 -8.530 ;
        RECT 97.770 -8.230 98.920 -8.150 ;
        RECT 105.210 -8.150 105.660 -8.050 ;
        RECT 111.970 -5.100 112.420 -5.000 ;
        RECT 118.710 -5.000 119.860 -4.920 ;
        RECT 124.770 -4.620 125.920 -4.540 ;
        RECT 132.210 -4.540 132.660 -4.440 ;
        RECT 138.970 -1.490 139.420 -1.390 ;
        RECT 145.710 -1.390 146.860 -1.310 ;
        RECT 151.770 -1.010 152.920 -0.930 ;
        RECT 159.210 -0.930 159.660 -0.830 ;
        RECT 165.970 2.120 166.420 2.220 ;
        RECT 172.710 2.220 173.860 2.300 ;
        RECT 178.770 2.600 179.920 2.680 ;
        RECT 186.210 2.680 186.660 2.780 ;
        RECT 192.970 5.730 193.420 5.830 ;
        RECT 199.710 5.830 200.860 5.910 ;
        RECT 205.770 6.210 206.920 6.290 ;
        RECT 213.210 6.290 213.660 6.390 ;
        RECT 207.170 6.210 207.580 6.270 ;
        RECT 205.770 5.910 207.580 6.210 ;
        RECT 205.770 5.830 206.920 5.910 ;
        RECT 207.170 5.850 207.580 5.910 ;
        RECT 212.550 6.210 212.960 6.270 ;
        RECT 213.210 6.210 214.360 6.290 ;
        RECT 212.550 5.910 214.360 6.210 ;
        RECT 212.550 5.850 212.960 5.910 ;
        RECT 199.710 5.730 200.160 5.830 ;
        RECT 192.970 4.580 193.410 5.730 ;
        RECT 199.720 4.580 200.160 5.730 ;
        RECT 192.970 3.930 194.120 4.580 ;
        RECT 199.010 3.930 200.160 4.580 ;
        RECT 192.970 2.780 193.410 3.930 ;
        RECT 199.720 2.780 200.160 3.930 ;
        RECT 192.970 2.680 193.420 2.780 ;
        RECT 180.170 2.600 180.580 2.660 ;
        RECT 178.770 2.300 180.580 2.600 ;
        RECT 178.770 2.220 179.920 2.300 ;
        RECT 180.170 2.240 180.580 2.300 ;
        RECT 185.550 2.600 185.960 2.660 ;
        RECT 186.210 2.600 187.360 2.680 ;
        RECT 185.550 2.300 187.360 2.600 ;
        RECT 185.550 2.240 185.960 2.300 ;
        RECT 172.710 2.120 173.160 2.220 ;
        RECT 165.970 0.970 166.410 2.120 ;
        RECT 172.720 0.970 173.160 2.120 ;
        RECT 165.970 0.320 167.120 0.970 ;
        RECT 172.010 0.320 173.160 0.970 ;
        RECT 165.970 -0.830 166.410 0.320 ;
        RECT 172.720 -0.830 173.160 0.320 ;
        RECT 165.970 -0.930 166.420 -0.830 ;
        RECT 153.170 -1.010 153.580 -0.950 ;
        RECT 151.770 -1.310 153.580 -1.010 ;
        RECT 151.770 -1.390 152.920 -1.310 ;
        RECT 153.170 -1.370 153.580 -1.310 ;
        RECT 158.550 -1.010 158.960 -0.950 ;
        RECT 159.210 -1.010 160.360 -0.930 ;
        RECT 158.550 -1.310 160.360 -1.010 ;
        RECT 158.550 -1.370 158.960 -1.310 ;
        RECT 145.710 -1.490 146.160 -1.390 ;
        RECT 138.970 -2.640 139.410 -1.490 ;
        RECT 145.720 -2.640 146.160 -1.490 ;
        RECT 138.970 -3.290 140.120 -2.640 ;
        RECT 145.010 -3.290 146.160 -2.640 ;
        RECT 138.970 -4.440 139.410 -3.290 ;
        RECT 145.720 -4.440 146.160 -3.290 ;
        RECT 138.970 -4.540 139.420 -4.440 ;
        RECT 126.170 -4.620 126.580 -4.560 ;
        RECT 124.770 -4.920 126.580 -4.620 ;
        RECT 124.770 -5.000 125.920 -4.920 ;
        RECT 126.170 -4.980 126.580 -4.920 ;
        RECT 131.550 -4.620 131.960 -4.560 ;
        RECT 132.210 -4.620 133.360 -4.540 ;
        RECT 131.550 -4.920 133.360 -4.620 ;
        RECT 131.550 -4.980 131.960 -4.920 ;
        RECT 118.710 -5.100 119.160 -5.000 ;
        RECT 111.970 -6.250 112.410 -5.100 ;
        RECT 118.720 -6.250 119.160 -5.100 ;
        RECT 111.970 -6.900 113.120 -6.250 ;
        RECT 118.010 -6.900 119.160 -6.250 ;
        RECT 111.970 -8.050 112.410 -6.900 ;
        RECT 118.720 -8.050 119.160 -6.900 ;
        RECT 111.970 -8.150 112.420 -8.050 ;
        RECT 99.170 -8.230 99.580 -8.170 ;
        RECT 97.770 -8.530 99.580 -8.230 ;
        RECT 97.770 -8.610 98.920 -8.530 ;
        RECT 99.170 -8.590 99.580 -8.530 ;
        RECT 104.550 -8.230 104.960 -8.170 ;
        RECT 105.210 -8.230 106.360 -8.150 ;
        RECT 104.550 -8.530 106.360 -8.230 ;
        RECT 104.550 -8.590 104.960 -8.530 ;
        RECT 91.710 -8.710 92.160 -8.610 ;
        RECT 84.970 -9.860 85.410 -8.710 ;
        RECT 91.720 -9.860 92.160 -8.710 ;
        RECT 84.970 -10.510 86.120 -9.860 ;
        RECT 91.010 -10.510 92.160 -9.860 ;
        RECT 84.970 -11.660 85.410 -10.510 ;
        RECT 91.720 -11.660 92.160 -10.510 ;
        RECT 84.970 -11.760 85.420 -11.660 ;
        RECT 72.170 -11.840 72.580 -11.780 ;
        RECT 70.770 -12.140 72.580 -11.840 ;
        RECT 70.770 -12.220 71.920 -12.140 ;
        RECT 72.170 -12.200 72.580 -12.140 ;
        RECT 77.550 -11.840 77.960 -11.780 ;
        RECT 78.210 -11.840 79.360 -11.760 ;
        RECT 77.550 -12.140 79.360 -11.840 ;
        RECT 77.550 -12.200 77.960 -12.140 ;
        RECT 64.710 -12.320 65.160 -12.220 ;
        RECT 57.970 -13.470 58.410 -12.320 ;
        RECT 64.720 -13.470 65.160 -12.320 ;
        RECT 57.970 -14.120 59.120 -13.470 ;
        RECT 64.010 -14.120 65.160 -13.470 ;
        RECT 57.970 -15.270 58.410 -14.120 ;
        RECT 64.720 -15.270 65.160 -14.120 ;
        RECT 57.970 -15.370 58.420 -15.270 ;
        RECT 45.170 -15.450 45.580 -15.390 ;
        RECT 43.770 -15.750 45.580 -15.450 ;
        RECT 43.770 -15.830 44.920 -15.750 ;
        RECT 45.170 -15.810 45.580 -15.750 ;
        RECT 50.550 -15.450 50.960 -15.390 ;
        RECT 51.210 -15.450 52.360 -15.370 ;
        RECT 50.550 -15.750 52.360 -15.450 ;
        RECT 50.550 -15.810 50.960 -15.750 ;
        RECT 37.710 -15.930 38.160 -15.830 ;
        RECT 30.970 -17.080 31.410 -15.930 ;
        RECT 37.720 -17.080 38.160 -15.930 ;
        RECT 30.970 -17.730 32.120 -17.080 ;
        RECT 37.010 -17.730 38.160 -17.080 ;
        RECT 30.970 -18.880 31.410 -17.730 ;
        RECT 37.720 -18.880 38.160 -17.730 ;
        RECT 30.970 -18.980 31.420 -18.880 ;
        RECT 18.170 -19.060 18.580 -19.000 ;
        RECT 16.770 -19.360 18.580 -19.060 ;
        RECT 16.770 -19.440 17.920 -19.360 ;
        RECT 18.170 -19.420 18.580 -19.360 ;
        RECT 23.550 -19.060 23.960 -19.000 ;
        RECT 24.210 -19.060 25.360 -18.980 ;
        RECT 23.550 -19.360 25.360 -19.060 ;
        RECT 23.550 -19.420 23.960 -19.360 ;
        RECT 10.710 -19.540 11.160 -19.440 ;
        RECT 3.970 -20.690 4.410 -19.540 ;
        RECT 10.720 -20.690 11.160 -19.540 ;
        RECT 3.970 -21.340 5.120 -20.690 ;
        RECT 10.010 -21.340 11.160 -20.690 ;
        RECT 3.970 -22.490 4.410 -21.340 ;
        RECT 10.720 -22.490 11.160 -21.340 ;
        RECT 3.970 -22.590 4.420 -22.490 ;
        RECT 3.270 -22.670 4.420 -22.590 ;
        RECT 10.710 -22.590 11.160 -22.490 ;
        RECT 17.470 -19.540 17.920 -19.440 ;
        RECT 24.210 -19.440 25.360 -19.360 ;
        RECT 30.270 -19.060 31.420 -18.980 ;
        RECT 37.710 -18.980 38.160 -18.880 ;
        RECT 44.470 -15.930 44.920 -15.830 ;
        RECT 51.210 -15.830 52.360 -15.750 ;
        RECT 57.270 -15.450 58.420 -15.370 ;
        RECT 64.710 -15.370 65.160 -15.270 ;
        RECT 71.470 -12.320 71.920 -12.220 ;
        RECT 78.210 -12.220 79.360 -12.140 ;
        RECT 84.270 -11.840 85.420 -11.760 ;
        RECT 91.710 -11.760 92.160 -11.660 ;
        RECT 98.470 -8.710 98.920 -8.610 ;
        RECT 105.210 -8.610 106.360 -8.530 ;
        RECT 111.270 -8.230 112.420 -8.150 ;
        RECT 118.710 -8.150 119.160 -8.050 ;
        RECT 125.470 -5.100 125.920 -5.000 ;
        RECT 132.210 -5.000 133.360 -4.920 ;
        RECT 138.270 -4.620 139.420 -4.540 ;
        RECT 145.710 -4.540 146.160 -4.440 ;
        RECT 152.470 -1.490 152.920 -1.390 ;
        RECT 159.210 -1.390 160.360 -1.310 ;
        RECT 165.270 -1.010 166.420 -0.930 ;
        RECT 172.710 -0.930 173.160 -0.830 ;
        RECT 179.470 2.120 179.920 2.220 ;
        RECT 186.210 2.220 187.360 2.300 ;
        RECT 192.270 2.600 193.420 2.680 ;
        RECT 199.710 2.680 200.160 2.780 ;
        RECT 206.470 5.730 206.920 5.830 ;
        RECT 213.210 5.830 214.360 5.910 ;
        RECT 213.210 5.730 213.660 5.830 ;
        RECT 206.470 4.580 206.910 5.730 ;
        RECT 213.220 4.580 213.660 5.730 ;
        RECT 206.470 3.930 207.620 4.580 ;
        RECT 212.510 3.930 213.660 4.580 ;
        RECT 206.470 2.780 206.910 3.930 ;
        RECT 213.220 2.780 213.660 3.930 ;
        RECT 206.470 2.680 206.920 2.780 ;
        RECT 193.670 2.600 194.080 2.660 ;
        RECT 192.270 2.300 194.080 2.600 ;
        RECT 192.270 2.220 193.420 2.300 ;
        RECT 193.670 2.240 194.080 2.300 ;
        RECT 199.050 2.600 199.460 2.660 ;
        RECT 199.710 2.600 200.860 2.680 ;
        RECT 199.050 2.300 200.860 2.600 ;
        RECT 199.050 2.240 199.460 2.300 ;
        RECT 186.210 2.120 186.660 2.220 ;
        RECT 179.470 0.970 179.910 2.120 ;
        RECT 186.220 0.970 186.660 2.120 ;
        RECT 179.470 0.320 180.620 0.970 ;
        RECT 185.510 0.320 186.660 0.970 ;
        RECT 179.470 -0.830 179.910 0.320 ;
        RECT 186.220 -0.830 186.660 0.320 ;
        RECT 179.470 -0.930 179.920 -0.830 ;
        RECT 166.670 -1.010 167.080 -0.950 ;
        RECT 165.270 -1.310 167.080 -1.010 ;
        RECT 165.270 -1.390 166.420 -1.310 ;
        RECT 166.670 -1.370 167.080 -1.310 ;
        RECT 172.050 -1.010 172.460 -0.950 ;
        RECT 172.710 -1.010 173.860 -0.930 ;
        RECT 172.050 -1.310 173.860 -1.010 ;
        RECT 172.050 -1.370 172.460 -1.310 ;
        RECT 159.210 -1.490 159.660 -1.390 ;
        RECT 152.470 -2.640 152.910 -1.490 ;
        RECT 159.220 -2.640 159.660 -1.490 ;
        RECT 152.470 -3.290 153.620 -2.640 ;
        RECT 158.510 -3.290 159.660 -2.640 ;
        RECT 152.470 -4.440 152.910 -3.290 ;
        RECT 159.220 -4.440 159.660 -3.290 ;
        RECT 152.470 -4.540 152.920 -4.440 ;
        RECT 139.670 -4.620 140.080 -4.560 ;
        RECT 138.270 -4.920 140.080 -4.620 ;
        RECT 138.270 -5.000 139.420 -4.920 ;
        RECT 139.670 -4.980 140.080 -4.920 ;
        RECT 145.050 -4.620 145.460 -4.560 ;
        RECT 145.710 -4.620 146.860 -4.540 ;
        RECT 145.050 -4.920 146.860 -4.620 ;
        RECT 145.050 -4.980 145.460 -4.920 ;
        RECT 132.210 -5.100 132.660 -5.000 ;
        RECT 125.470 -6.250 125.910 -5.100 ;
        RECT 132.220 -6.250 132.660 -5.100 ;
        RECT 125.470 -6.900 126.620 -6.250 ;
        RECT 131.510 -6.900 132.660 -6.250 ;
        RECT 125.470 -8.050 125.910 -6.900 ;
        RECT 132.220 -8.050 132.660 -6.900 ;
        RECT 125.470 -8.150 125.920 -8.050 ;
        RECT 112.670 -8.230 113.080 -8.170 ;
        RECT 111.270 -8.530 113.080 -8.230 ;
        RECT 111.270 -8.610 112.420 -8.530 ;
        RECT 112.670 -8.590 113.080 -8.530 ;
        RECT 118.050 -8.230 118.460 -8.170 ;
        RECT 118.710 -8.230 119.860 -8.150 ;
        RECT 118.050 -8.530 119.860 -8.230 ;
        RECT 118.050 -8.590 118.460 -8.530 ;
        RECT 105.210 -8.710 105.660 -8.610 ;
        RECT 98.470 -9.860 98.910 -8.710 ;
        RECT 105.220 -9.860 105.660 -8.710 ;
        RECT 98.470 -10.510 99.620 -9.860 ;
        RECT 104.510 -10.510 105.660 -9.860 ;
        RECT 98.470 -11.660 98.910 -10.510 ;
        RECT 105.220 -11.660 105.660 -10.510 ;
        RECT 98.470 -11.760 98.920 -11.660 ;
        RECT 85.670 -11.840 86.080 -11.780 ;
        RECT 84.270 -12.140 86.080 -11.840 ;
        RECT 84.270 -12.220 85.420 -12.140 ;
        RECT 85.670 -12.200 86.080 -12.140 ;
        RECT 91.050 -11.840 91.460 -11.780 ;
        RECT 91.710 -11.840 92.860 -11.760 ;
        RECT 91.050 -12.140 92.860 -11.840 ;
        RECT 91.050 -12.200 91.460 -12.140 ;
        RECT 78.210 -12.320 78.660 -12.220 ;
        RECT 71.470 -13.470 71.910 -12.320 ;
        RECT 78.220 -13.470 78.660 -12.320 ;
        RECT 71.470 -14.120 72.620 -13.470 ;
        RECT 77.510 -14.120 78.660 -13.470 ;
        RECT 71.470 -15.270 71.910 -14.120 ;
        RECT 78.220 -15.270 78.660 -14.120 ;
        RECT 71.470 -15.370 71.920 -15.270 ;
        RECT 58.670 -15.450 59.080 -15.390 ;
        RECT 57.270 -15.750 59.080 -15.450 ;
        RECT 57.270 -15.830 58.420 -15.750 ;
        RECT 58.670 -15.810 59.080 -15.750 ;
        RECT 64.050 -15.450 64.460 -15.390 ;
        RECT 64.710 -15.450 65.860 -15.370 ;
        RECT 64.050 -15.750 65.860 -15.450 ;
        RECT 64.050 -15.810 64.460 -15.750 ;
        RECT 51.210 -15.930 51.660 -15.830 ;
        RECT 44.470 -17.080 44.910 -15.930 ;
        RECT 51.220 -17.080 51.660 -15.930 ;
        RECT 44.470 -17.730 45.620 -17.080 ;
        RECT 50.510 -17.730 51.660 -17.080 ;
        RECT 44.470 -18.880 44.910 -17.730 ;
        RECT 51.220 -18.880 51.660 -17.730 ;
        RECT 44.470 -18.980 44.920 -18.880 ;
        RECT 31.670 -19.060 32.080 -19.000 ;
        RECT 30.270 -19.360 32.080 -19.060 ;
        RECT 30.270 -19.440 31.420 -19.360 ;
        RECT 31.670 -19.420 32.080 -19.360 ;
        RECT 37.050 -19.060 37.460 -19.000 ;
        RECT 37.710 -19.060 38.860 -18.980 ;
        RECT 37.050 -19.360 38.860 -19.060 ;
        RECT 37.050 -19.420 37.460 -19.360 ;
        RECT 24.210 -19.540 24.660 -19.440 ;
        RECT 17.470 -20.690 17.910 -19.540 ;
        RECT 24.220 -20.690 24.660 -19.540 ;
        RECT 17.470 -21.340 18.620 -20.690 ;
        RECT 23.510 -21.340 24.660 -20.690 ;
        RECT 17.470 -22.490 17.910 -21.340 ;
        RECT 24.220 -22.490 24.660 -21.340 ;
        RECT 17.470 -22.590 17.920 -22.490 ;
        RECT 4.670 -22.670 5.080 -22.610 ;
        RECT 3.270 -22.970 5.080 -22.670 ;
        RECT 3.270 -23.050 4.420 -22.970 ;
        RECT 4.670 -23.030 5.080 -22.970 ;
        RECT 10.050 -22.670 10.460 -22.610 ;
        RECT 10.710 -22.670 11.860 -22.590 ;
        RECT 10.050 -22.970 11.860 -22.670 ;
        RECT 10.050 -23.030 10.460 -22.970 ;
        RECT 3.970 -23.150 4.420 -23.050 ;
        RECT 10.710 -23.050 11.860 -22.970 ;
        RECT 16.770 -22.670 17.920 -22.590 ;
        RECT 24.210 -22.590 24.660 -22.490 ;
        RECT 30.970 -19.540 31.420 -19.440 ;
        RECT 37.710 -19.440 38.860 -19.360 ;
        RECT 43.770 -19.060 44.920 -18.980 ;
        RECT 51.210 -18.980 51.660 -18.880 ;
        RECT 57.970 -15.930 58.420 -15.830 ;
        RECT 64.710 -15.830 65.860 -15.750 ;
        RECT 70.770 -15.450 71.920 -15.370 ;
        RECT 78.210 -15.370 78.660 -15.270 ;
        RECT 84.970 -12.320 85.420 -12.220 ;
        RECT 91.710 -12.220 92.860 -12.140 ;
        RECT 97.770 -11.840 98.920 -11.760 ;
        RECT 105.210 -11.760 105.660 -11.660 ;
        RECT 111.970 -8.710 112.420 -8.610 ;
        RECT 118.710 -8.610 119.860 -8.530 ;
        RECT 124.770 -8.230 125.920 -8.150 ;
        RECT 132.210 -8.150 132.660 -8.050 ;
        RECT 138.970 -5.100 139.420 -5.000 ;
        RECT 145.710 -5.000 146.860 -4.920 ;
        RECT 151.770 -4.620 152.920 -4.540 ;
        RECT 159.210 -4.540 159.660 -4.440 ;
        RECT 165.970 -1.490 166.420 -1.390 ;
        RECT 172.710 -1.390 173.860 -1.310 ;
        RECT 178.770 -1.010 179.920 -0.930 ;
        RECT 186.210 -0.930 186.660 -0.830 ;
        RECT 192.970 2.120 193.420 2.220 ;
        RECT 199.710 2.220 200.860 2.300 ;
        RECT 205.770 2.600 206.920 2.680 ;
        RECT 213.210 2.680 213.660 2.780 ;
        RECT 207.170 2.600 207.580 2.660 ;
        RECT 205.770 2.300 207.580 2.600 ;
        RECT 205.770 2.220 206.920 2.300 ;
        RECT 207.170 2.240 207.580 2.300 ;
        RECT 212.550 2.600 212.960 2.660 ;
        RECT 213.210 2.600 214.360 2.680 ;
        RECT 212.550 2.300 214.360 2.600 ;
        RECT 212.550 2.240 212.960 2.300 ;
        RECT 199.710 2.120 200.160 2.220 ;
        RECT 192.970 0.970 193.410 2.120 ;
        RECT 199.720 0.970 200.160 2.120 ;
        RECT 192.970 0.320 194.120 0.970 ;
        RECT 199.010 0.320 200.160 0.970 ;
        RECT 192.970 -0.830 193.410 0.320 ;
        RECT 199.720 -0.830 200.160 0.320 ;
        RECT 192.970 -0.930 193.420 -0.830 ;
        RECT 180.170 -1.010 180.580 -0.950 ;
        RECT 178.770 -1.310 180.580 -1.010 ;
        RECT 178.770 -1.390 179.920 -1.310 ;
        RECT 180.170 -1.370 180.580 -1.310 ;
        RECT 185.550 -1.010 185.960 -0.950 ;
        RECT 186.210 -1.010 187.360 -0.930 ;
        RECT 185.550 -1.310 187.360 -1.010 ;
        RECT 185.550 -1.370 185.960 -1.310 ;
        RECT 172.710 -1.490 173.160 -1.390 ;
        RECT 165.970 -2.640 166.410 -1.490 ;
        RECT 172.720 -2.640 173.160 -1.490 ;
        RECT 165.970 -3.290 167.120 -2.640 ;
        RECT 172.010 -3.290 173.160 -2.640 ;
        RECT 165.970 -4.440 166.410 -3.290 ;
        RECT 172.720 -4.440 173.160 -3.290 ;
        RECT 165.970 -4.540 166.420 -4.440 ;
        RECT 153.170 -4.620 153.580 -4.560 ;
        RECT 151.770 -4.920 153.580 -4.620 ;
        RECT 151.770 -5.000 152.920 -4.920 ;
        RECT 153.170 -4.980 153.580 -4.920 ;
        RECT 158.550 -4.620 158.960 -4.560 ;
        RECT 159.210 -4.620 160.360 -4.540 ;
        RECT 158.550 -4.920 160.360 -4.620 ;
        RECT 158.550 -4.980 158.960 -4.920 ;
        RECT 145.710 -5.100 146.160 -5.000 ;
        RECT 138.970 -6.250 139.410 -5.100 ;
        RECT 145.720 -6.250 146.160 -5.100 ;
        RECT 138.970 -6.900 140.120 -6.250 ;
        RECT 145.010 -6.900 146.160 -6.250 ;
        RECT 138.970 -8.050 139.410 -6.900 ;
        RECT 145.720 -8.050 146.160 -6.900 ;
        RECT 138.970 -8.150 139.420 -8.050 ;
        RECT 126.170 -8.230 126.580 -8.170 ;
        RECT 124.770 -8.530 126.580 -8.230 ;
        RECT 124.770 -8.610 125.920 -8.530 ;
        RECT 126.170 -8.590 126.580 -8.530 ;
        RECT 131.550 -8.230 131.960 -8.170 ;
        RECT 132.210 -8.230 133.360 -8.150 ;
        RECT 131.550 -8.530 133.360 -8.230 ;
        RECT 131.550 -8.590 131.960 -8.530 ;
        RECT 118.710 -8.710 119.160 -8.610 ;
        RECT 111.970 -9.860 112.410 -8.710 ;
        RECT 118.720 -9.860 119.160 -8.710 ;
        RECT 111.970 -10.510 113.120 -9.860 ;
        RECT 118.010 -10.510 119.160 -9.860 ;
        RECT 111.970 -11.660 112.410 -10.510 ;
        RECT 118.720 -11.660 119.160 -10.510 ;
        RECT 111.970 -11.760 112.420 -11.660 ;
        RECT 99.170 -11.840 99.580 -11.780 ;
        RECT 97.770 -12.140 99.580 -11.840 ;
        RECT 97.770 -12.220 98.920 -12.140 ;
        RECT 99.170 -12.200 99.580 -12.140 ;
        RECT 104.550 -11.840 104.960 -11.780 ;
        RECT 105.210 -11.840 106.360 -11.760 ;
        RECT 104.550 -12.140 106.360 -11.840 ;
        RECT 104.550 -12.200 104.960 -12.140 ;
        RECT 91.710 -12.320 92.160 -12.220 ;
        RECT 84.970 -13.470 85.410 -12.320 ;
        RECT 91.720 -13.470 92.160 -12.320 ;
        RECT 84.970 -14.120 86.120 -13.470 ;
        RECT 91.010 -14.120 92.160 -13.470 ;
        RECT 84.970 -15.270 85.410 -14.120 ;
        RECT 91.720 -15.270 92.160 -14.120 ;
        RECT 84.970 -15.370 85.420 -15.270 ;
        RECT 72.170 -15.450 72.580 -15.390 ;
        RECT 70.770 -15.750 72.580 -15.450 ;
        RECT 70.770 -15.830 71.920 -15.750 ;
        RECT 72.170 -15.810 72.580 -15.750 ;
        RECT 77.550 -15.450 77.960 -15.390 ;
        RECT 78.210 -15.450 79.360 -15.370 ;
        RECT 77.550 -15.750 79.360 -15.450 ;
        RECT 77.550 -15.810 77.960 -15.750 ;
        RECT 64.710 -15.930 65.160 -15.830 ;
        RECT 57.970 -17.080 58.410 -15.930 ;
        RECT 64.720 -17.080 65.160 -15.930 ;
        RECT 57.970 -17.730 59.120 -17.080 ;
        RECT 64.010 -17.730 65.160 -17.080 ;
        RECT 57.970 -18.880 58.410 -17.730 ;
        RECT 64.720 -18.880 65.160 -17.730 ;
        RECT 57.970 -18.980 58.420 -18.880 ;
        RECT 45.170 -19.060 45.580 -19.000 ;
        RECT 43.770 -19.360 45.580 -19.060 ;
        RECT 43.770 -19.440 44.920 -19.360 ;
        RECT 45.170 -19.420 45.580 -19.360 ;
        RECT 50.550 -19.060 50.960 -19.000 ;
        RECT 51.210 -19.060 52.360 -18.980 ;
        RECT 50.550 -19.360 52.360 -19.060 ;
        RECT 50.550 -19.420 50.960 -19.360 ;
        RECT 37.710 -19.540 38.160 -19.440 ;
        RECT 30.970 -20.690 31.410 -19.540 ;
        RECT 37.720 -20.690 38.160 -19.540 ;
        RECT 30.970 -21.340 32.120 -20.690 ;
        RECT 37.010 -21.340 38.160 -20.690 ;
        RECT 30.970 -22.490 31.410 -21.340 ;
        RECT 37.720 -22.490 38.160 -21.340 ;
        RECT 30.970 -22.590 31.420 -22.490 ;
        RECT 18.170 -22.670 18.580 -22.610 ;
        RECT 16.770 -22.970 18.580 -22.670 ;
        RECT 16.770 -23.050 17.920 -22.970 ;
        RECT 18.170 -23.030 18.580 -22.970 ;
        RECT 23.550 -22.670 23.960 -22.610 ;
        RECT 24.210 -22.670 25.360 -22.590 ;
        RECT 23.550 -22.970 25.360 -22.670 ;
        RECT 23.550 -23.030 23.960 -22.970 ;
        RECT 10.710 -23.150 11.160 -23.050 ;
        RECT 3.970 -24.300 4.410 -23.150 ;
        RECT 10.720 -24.300 11.160 -23.150 ;
        RECT 3.970 -24.950 5.120 -24.300 ;
        RECT 10.010 -24.950 11.160 -24.300 ;
        RECT 3.970 -26.100 4.410 -24.950 ;
        RECT 10.720 -26.100 11.160 -24.950 ;
        RECT 3.970 -26.200 4.420 -26.100 ;
        RECT 3.270 -26.280 4.420 -26.200 ;
        RECT 10.710 -26.200 11.160 -26.100 ;
        RECT 17.470 -23.150 17.920 -23.050 ;
        RECT 24.210 -23.050 25.360 -22.970 ;
        RECT 30.270 -22.670 31.420 -22.590 ;
        RECT 37.710 -22.590 38.160 -22.490 ;
        RECT 44.470 -19.540 44.920 -19.440 ;
        RECT 51.210 -19.440 52.360 -19.360 ;
        RECT 57.270 -19.060 58.420 -18.980 ;
        RECT 64.710 -18.980 65.160 -18.880 ;
        RECT 71.470 -15.930 71.920 -15.830 ;
        RECT 78.210 -15.830 79.360 -15.750 ;
        RECT 84.270 -15.450 85.420 -15.370 ;
        RECT 91.710 -15.370 92.160 -15.270 ;
        RECT 98.470 -12.320 98.920 -12.220 ;
        RECT 105.210 -12.220 106.360 -12.140 ;
        RECT 111.270 -11.840 112.420 -11.760 ;
        RECT 118.710 -11.760 119.160 -11.660 ;
        RECT 125.470 -8.710 125.920 -8.610 ;
        RECT 132.210 -8.610 133.360 -8.530 ;
        RECT 138.270 -8.230 139.420 -8.150 ;
        RECT 145.710 -8.150 146.160 -8.050 ;
        RECT 152.470 -5.100 152.920 -5.000 ;
        RECT 159.210 -5.000 160.360 -4.920 ;
        RECT 165.270 -4.620 166.420 -4.540 ;
        RECT 172.710 -4.540 173.160 -4.440 ;
        RECT 179.470 -1.490 179.920 -1.390 ;
        RECT 186.210 -1.390 187.360 -1.310 ;
        RECT 192.270 -1.010 193.420 -0.930 ;
        RECT 199.710 -0.930 200.160 -0.830 ;
        RECT 206.470 2.120 206.920 2.220 ;
        RECT 213.210 2.220 214.360 2.300 ;
        RECT 213.210 2.120 213.660 2.220 ;
        RECT 206.470 0.970 206.910 2.120 ;
        RECT 213.220 0.970 213.660 2.120 ;
        RECT 206.470 0.320 207.620 0.970 ;
        RECT 212.510 0.320 213.660 0.970 ;
        RECT 206.470 -0.830 206.910 0.320 ;
        RECT 213.220 -0.830 213.660 0.320 ;
        RECT 206.470 -0.930 206.920 -0.830 ;
        RECT 193.670 -1.010 194.080 -0.950 ;
        RECT 192.270 -1.310 194.080 -1.010 ;
        RECT 192.270 -1.390 193.420 -1.310 ;
        RECT 193.670 -1.370 194.080 -1.310 ;
        RECT 199.050 -1.010 199.460 -0.950 ;
        RECT 199.710 -1.010 200.860 -0.930 ;
        RECT 199.050 -1.310 200.860 -1.010 ;
        RECT 199.050 -1.370 199.460 -1.310 ;
        RECT 186.210 -1.490 186.660 -1.390 ;
        RECT 179.470 -2.640 179.910 -1.490 ;
        RECT 186.220 -2.640 186.660 -1.490 ;
        RECT 179.470 -3.290 180.620 -2.640 ;
        RECT 185.510 -3.290 186.660 -2.640 ;
        RECT 179.470 -4.440 179.910 -3.290 ;
        RECT 186.220 -4.440 186.660 -3.290 ;
        RECT 179.470 -4.540 179.920 -4.440 ;
        RECT 166.670 -4.620 167.080 -4.560 ;
        RECT 165.270 -4.920 167.080 -4.620 ;
        RECT 165.270 -5.000 166.420 -4.920 ;
        RECT 166.670 -4.980 167.080 -4.920 ;
        RECT 172.050 -4.620 172.460 -4.560 ;
        RECT 172.710 -4.620 173.860 -4.540 ;
        RECT 172.050 -4.920 173.860 -4.620 ;
        RECT 172.050 -4.980 172.460 -4.920 ;
        RECT 159.210 -5.100 159.660 -5.000 ;
        RECT 152.470 -6.250 152.910 -5.100 ;
        RECT 159.220 -6.250 159.660 -5.100 ;
        RECT 152.470 -6.900 153.620 -6.250 ;
        RECT 158.510 -6.900 159.660 -6.250 ;
        RECT 152.470 -8.050 152.910 -6.900 ;
        RECT 159.220 -8.050 159.660 -6.900 ;
        RECT 152.470 -8.150 152.920 -8.050 ;
        RECT 139.670 -8.230 140.080 -8.170 ;
        RECT 138.270 -8.530 140.080 -8.230 ;
        RECT 138.270 -8.610 139.420 -8.530 ;
        RECT 139.670 -8.590 140.080 -8.530 ;
        RECT 145.050 -8.230 145.460 -8.170 ;
        RECT 145.710 -8.230 146.860 -8.150 ;
        RECT 145.050 -8.530 146.860 -8.230 ;
        RECT 145.050 -8.590 145.460 -8.530 ;
        RECT 132.210 -8.710 132.660 -8.610 ;
        RECT 125.470 -9.860 125.910 -8.710 ;
        RECT 132.220 -9.860 132.660 -8.710 ;
        RECT 125.470 -10.510 126.620 -9.860 ;
        RECT 131.510 -10.510 132.660 -9.860 ;
        RECT 125.470 -11.660 125.910 -10.510 ;
        RECT 132.220 -11.660 132.660 -10.510 ;
        RECT 125.470 -11.760 125.920 -11.660 ;
        RECT 112.670 -11.840 113.080 -11.780 ;
        RECT 111.270 -12.140 113.080 -11.840 ;
        RECT 111.270 -12.220 112.420 -12.140 ;
        RECT 112.670 -12.200 113.080 -12.140 ;
        RECT 118.050 -11.840 118.460 -11.780 ;
        RECT 118.710 -11.840 119.860 -11.760 ;
        RECT 118.050 -12.140 119.860 -11.840 ;
        RECT 118.050 -12.200 118.460 -12.140 ;
        RECT 105.210 -12.320 105.660 -12.220 ;
        RECT 98.470 -13.470 98.910 -12.320 ;
        RECT 105.220 -13.470 105.660 -12.320 ;
        RECT 98.470 -14.120 99.620 -13.470 ;
        RECT 104.510 -14.120 105.660 -13.470 ;
        RECT 98.470 -15.270 98.910 -14.120 ;
        RECT 105.220 -15.270 105.660 -14.120 ;
        RECT 98.470 -15.370 98.920 -15.270 ;
        RECT 85.670 -15.450 86.080 -15.390 ;
        RECT 84.270 -15.750 86.080 -15.450 ;
        RECT 84.270 -15.830 85.420 -15.750 ;
        RECT 85.670 -15.810 86.080 -15.750 ;
        RECT 91.050 -15.450 91.460 -15.390 ;
        RECT 91.710 -15.450 92.860 -15.370 ;
        RECT 91.050 -15.750 92.860 -15.450 ;
        RECT 91.050 -15.810 91.460 -15.750 ;
        RECT 78.210 -15.930 78.660 -15.830 ;
        RECT 71.470 -17.080 71.910 -15.930 ;
        RECT 78.220 -17.080 78.660 -15.930 ;
        RECT 71.470 -17.730 72.620 -17.080 ;
        RECT 77.510 -17.730 78.660 -17.080 ;
        RECT 71.470 -18.880 71.910 -17.730 ;
        RECT 78.220 -18.880 78.660 -17.730 ;
        RECT 71.470 -18.980 71.920 -18.880 ;
        RECT 58.670 -19.060 59.080 -19.000 ;
        RECT 57.270 -19.360 59.080 -19.060 ;
        RECT 57.270 -19.440 58.420 -19.360 ;
        RECT 58.670 -19.420 59.080 -19.360 ;
        RECT 64.050 -19.060 64.460 -19.000 ;
        RECT 64.710 -19.060 65.860 -18.980 ;
        RECT 64.050 -19.360 65.860 -19.060 ;
        RECT 64.050 -19.420 64.460 -19.360 ;
        RECT 51.210 -19.540 51.660 -19.440 ;
        RECT 44.470 -20.690 44.910 -19.540 ;
        RECT 51.220 -20.690 51.660 -19.540 ;
        RECT 44.470 -21.340 45.620 -20.690 ;
        RECT 50.510 -21.340 51.660 -20.690 ;
        RECT 44.470 -22.490 44.910 -21.340 ;
        RECT 51.220 -22.490 51.660 -21.340 ;
        RECT 44.470 -22.590 44.920 -22.490 ;
        RECT 31.670 -22.670 32.080 -22.610 ;
        RECT 30.270 -22.970 32.080 -22.670 ;
        RECT 30.270 -23.050 31.420 -22.970 ;
        RECT 31.670 -23.030 32.080 -22.970 ;
        RECT 37.050 -22.670 37.460 -22.610 ;
        RECT 37.710 -22.670 38.860 -22.590 ;
        RECT 37.050 -22.970 38.860 -22.670 ;
        RECT 37.050 -23.030 37.460 -22.970 ;
        RECT 24.210 -23.150 24.660 -23.050 ;
        RECT 17.470 -24.300 17.910 -23.150 ;
        RECT 24.220 -24.300 24.660 -23.150 ;
        RECT 17.470 -24.950 18.620 -24.300 ;
        RECT 23.510 -24.950 24.660 -24.300 ;
        RECT 17.470 -26.100 17.910 -24.950 ;
        RECT 24.220 -26.100 24.660 -24.950 ;
        RECT 17.470 -26.200 17.920 -26.100 ;
        RECT 4.670 -26.280 5.080 -26.220 ;
        RECT 3.270 -26.580 5.080 -26.280 ;
        RECT 3.270 -26.660 4.420 -26.580 ;
        RECT 4.670 -26.640 5.080 -26.580 ;
        RECT 10.050 -26.280 10.460 -26.220 ;
        RECT 10.710 -26.280 11.860 -26.200 ;
        RECT 10.050 -26.580 11.860 -26.280 ;
        RECT 10.050 -26.640 10.460 -26.580 ;
        RECT 3.970 -26.760 4.420 -26.660 ;
        RECT 10.710 -26.660 11.860 -26.580 ;
        RECT 16.770 -26.280 17.920 -26.200 ;
        RECT 24.210 -26.200 24.660 -26.100 ;
        RECT 30.970 -23.150 31.420 -23.050 ;
        RECT 37.710 -23.050 38.860 -22.970 ;
        RECT 43.770 -22.670 44.920 -22.590 ;
        RECT 51.210 -22.590 51.660 -22.490 ;
        RECT 57.970 -19.540 58.420 -19.440 ;
        RECT 64.710 -19.440 65.860 -19.360 ;
        RECT 70.770 -19.060 71.920 -18.980 ;
        RECT 78.210 -18.980 78.660 -18.880 ;
        RECT 84.970 -15.930 85.420 -15.830 ;
        RECT 91.710 -15.830 92.860 -15.750 ;
        RECT 97.770 -15.450 98.920 -15.370 ;
        RECT 105.210 -15.370 105.660 -15.270 ;
        RECT 111.970 -12.320 112.420 -12.220 ;
        RECT 118.710 -12.220 119.860 -12.140 ;
        RECT 124.770 -11.840 125.920 -11.760 ;
        RECT 132.210 -11.760 132.660 -11.660 ;
        RECT 138.970 -8.710 139.420 -8.610 ;
        RECT 145.710 -8.610 146.860 -8.530 ;
        RECT 151.770 -8.230 152.920 -8.150 ;
        RECT 159.210 -8.150 159.660 -8.050 ;
        RECT 165.970 -5.100 166.420 -5.000 ;
        RECT 172.710 -5.000 173.860 -4.920 ;
        RECT 178.770 -4.620 179.920 -4.540 ;
        RECT 186.210 -4.540 186.660 -4.440 ;
        RECT 192.970 -1.490 193.420 -1.390 ;
        RECT 199.710 -1.390 200.860 -1.310 ;
        RECT 205.770 -1.010 206.920 -0.930 ;
        RECT 213.210 -0.930 213.660 -0.830 ;
        RECT 207.170 -1.010 207.580 -0.950 ;
        RECT 205.770 -1.310 207.580 -1.010 ;
        RECT 205.770 -1.390 206.920 -1.310 ;
        RECT 207.170 -1.370 207.580 -1.310 ;
        RECT 212.550 -1.010 212.960 -0.950 ;
        RECT 213.210 -1.010 214.360 -0.930 ;
        RECT 212.550 -1.310 214.360 -1.010 ;
        RECT 212.550 -1.370 212.960 -1.310 ;
        RECT 199.710 -1.490 200.160 -1.390 ;
        RECT 192.970 -2.640 193.410 -1.490 ;
        RECT 199.720 -2.640 200.160 -1.490 ;
        RECT 192.970 -3.290 194.120 -2.640 ;
        RECT 199.010 -3.290 200.160 -2.640 ;
        RECT 192.970 -4.440 193.410 -3.290 ;
        RECT 199.720 -4.440 200.160 -3.290 ;
        RECT 192.970 -4.540 193.420 -4.440 ;
        RECT 180.170 -4.620 180.580 -4.560 ;
        RECT 178.770 -4.920 180.580 -4.620 ;
        RECT 178.770 -5.000 179.920 -4.920 ;
        RECT 180.170 -4.980 180.580 -4.920 ;
        RECT 185.550 -4.620 185.960 -4.560 ;
        RECT 186.210 -4.620 187.360 -4.540 ;
        RECT 185.550 -4.920 187.360 -4.620 ;
        RECT 185.550 -4.980 185.960 -4.920 ;
        RECT 172.710 -5.100 173.160 -5.000 ;
        RECT 165.970 -6.250 166.410 -5.100 ;
        RECT 172.720 -6.250 173.160 -5.100 ;
        RECT 165.970 -6.900 167.120 -6.250 ;
        RECT 172.010 -6.900 173.160 -6.250 ;
        RECT 165.970 -8.050 166.410 -6.900 ;
        RECT 172.720 -8.050 173.160 -6.900 ;
        RECT 165.970 -8.150 166.420 -8.050 ;
        RECT 153.170 -8.230 153.580 -8.170 ;
        RECT 151.770 -8.530 153.580 -8.230 ;
        RECT 151.770 -8.610 152.920 -8.530 ;
        RECT 153.170 -8.590 153.580 -8.530 ;
        RECT 158.550 -8.230 158.960 -8.170 ;
        RECT 159.210 -8.230 160.360 -8.150 ;
        RECT 158.550 -8.530 160.360 -8.230 ;
        RECT 158.550 -8.590 158.960 -8.530 ;
        RECT 145.710 -8.710 146.160 -8.610 ;
        RECT 138.970 -9.860 139.410 -8.710 ;
        RECT 145.720 -9.860 146.160 -8.710 ;
        RECT 138.970 -10.510 140.120 -9.860 ;
        RECT 145.010 -10.510 146.160 -9.860 ;
        RECT 138.970 -11.660 139.410 -10.510 ;
        RECT 145.720 -11.660 146.160 -10.510 ;
        RECT 138.970 -11.760 139.420 -11.660 ;
        RECT 126.170 -11.840 126.580 -11.780 ;
        RECT 124.770 -12.140 126.580 -11.840 ;
        RECT 124.770 -12.220 125.920 -12.140 ;
        RECT 126.170 -12.200 126.580 -12.140 ;
        RECT 131.550 -11.840 131.960 -11.780 ;
        RECT 132.210 -11.840 133.360 -11.760 ;
        RECT 131.550 -12.140 133.360 -11.840 ;
        RECT 131.550 -12.200 131.960 -12.140 ;
        RECT 118.710 -12.320 119.160 -12.220 ;
        RECT 111.970 -13.470 112.410 -12.320 ;
        RECT 118.720 -13.470 119.160 -12.320 ;
        RECT 111.970 -14.120 113.120 -13.470 ;
        RECT 118.010 -14.120 119.160 -13.470 ;
        RECT 111.970 -15.270 112.410 -14.120 ;
        RECT 118.720 -15.270 119.160 -14.120 ;
        RECT 111.970 -15.370 112.420 -15.270 ;
        RECT 99.170 -15.450 99.580 -15.390 ;
        RECT 97.770 -15.750 99.580 -15.450 ;
        RECT 97.770 -15.830 98.920 -15.750 ;
        RECT 99.170 -15.810 99.580 -15.750 ;
        RECT 104.550 -15.450 104.960 -15.390 ;
        RECT 105.210 -15.450 106.360 -15.370 ;
        RECT 104.550 -15.750 106.360 -15.450 ;
        RECT 104.550 -15.810 104.960 -15.750 ;
        RECT 91.710 -15.930 92.160 -15.830 ;
        RECT 84.970 -17.080 85.410 -15.930 ;
        RECT 91.720 -17.080 92.160 -15.930 ;
        RECT 84.970 -17.730 86.120 -17.080 ;
        RECT 91.010 -17.730 92.160 -17.080 ;
        RECT 84.970 -18.880 85.410 -17.730 ;
        RECT 91.720 -18.880 92.160 -17.730 ;
        RECT 84.970 -18.980 85.420 -18.880 ;
        RECT 72.170 -19.060 72.580 -19.000 ;
        RECT 70.770 -19.360 72.580 -19.060 ;
        RECT 70.770 -19.440 71.920 -19.360 ;
        RECT 72.170 -19.420 72.580 -19.360 ;
        RECT 77.550 -19.060 77.960 -19.000 ;
        RECT 78.210 -19.060 79.360 -18.980 ;
        RECT 77.550 -19.360 79.360 -19.060 ;
        RECT 77.550 -19.420 77.960 -19.360 ;
        RECT 64.710 -19.540 65.160 -19.440 ;
        RECT 57.970 -20.690 58.410 -19.540 ;
        RECT 64.720 -20.690 65.160 -19.540 ;
        RECT 57.970 -21.340 59.120 -20.690 ;
        RECT 64.010 -21.340 65.160 -20.690 ;
        RECT 57.970 -22.490 58.410 -21.340 ;
        RECT 64.720 -22.490 65.160 -21.340 ;
        RECT 57.970 -22.590 58.420 -22.490 ;
        RECT 45.170 -22.670 45.580 -22.610 ;
        RECT 43.770 -22.970 45.580 -22.670 ;
        RECT 43.770 -23.050 44.920 -22.970 ;
        RECT 45.170 -23.030 45.580 -22.970 ;
        RECT 50.550 -22.670 50.960 -22.610 ;
        RECT 51.210 -22.670 52.360 -22.590 ;
        RECT 50.550 -22.970 52.360 -22.670 ;
        RECT 50.550 -23.030 50.960 -22.970 ;
        RECT 37.710 -23.150 38.160 -23.050 ;
        RECT 30.970 -24.300 31.410 -23.150 ;
        RECT 37.720 -24.300 38.160 -23.150 ;
        RECT 30.970 -24.950 32.120 -24.300 ;
        RECT 37.010 -24.950 38.160 -24.300 ;
        RECT 30.970 -26.100 31.410 -24.950 ;
        RECT 37.720 -26.100 38.160 -24.950 ;
        RECT 30.970 -26.200 31.420 -26.100 ;
        RECT 18.170 -26.280 18.580 -26.220 ;
        RECT 16.770 -26.580 18.580 -26.280 ;
        RECT 16.770 -26.660 17.920 -26.580 ;
        RECT 18.170 -26.640 18.580 -26.580 ;
        RECT 23.550 -26.280 23.960 -26.220 ;
        RECT 24.210 -26.280 25.360 -26.200 ;
        RECT 23.550 -26.580 25.360 -26.280 ;
        RECT 23.550 -26.640 23.960 -26.580 ;
        RECT 10.710 -26.760 11.160 -26.660 ;
        RECT 3.970 -27.910 4.410 -26.760 ;
        RECT 10.720 -27.910 11.160 -26.760 ;
        RECT 3.970 -28.560 5.120 -27.910 ;
        RECT 10.010 -28.560 11.160 -27.910 ;
        RECT 3.970 -29.710 4.410 -28.560 ;
        RECT 10.720 -29.710 11.160 -28.560 ;
        RECT 3.970 -29.810 4.420 -29.710 ;
        RECT 3.270 -29.890 4.420 -29.810 ;
        RECT 10.710 -29.810 11.160 -29.710 ;
        RECT 17.470 -26.760 17.920 -26.660 ;
        RECT 24.210 -26.660 25.360 -26.580 ;
        RECT 30.270 -26.280 31.420 -26.200 ;
        RECT 37.710 -26.200 38.160 -26.100 ;
        RECT 44.470 -23.150 44.920 -23.050 ;
        RECT 51.210 -23.050 52.360 -22.970 ;
        RECT 57.270 -22.670 58.420 -22.590 ;
        RECT 64.710 -22.590 65.160 -22.490 ;
        RECT 71.470 -19.540 71.920 -19.440 ;
        RECT 78.210 -19.440 79.360 -19.360 ;
        RECT 84.270 -19.060 85.420 -18.980 ;
        RECT 91.710 -18.980 92.160 -18.880 ;
        RECT 98.470 -15.930 98.920 -15.830 ;
        RECT 105.210 -15.830 106.360 -15.750 ;
        RECT 111.270 -15.450 112.420 -15.370 ;
        RECT 118.710 -15.370 119.160 -15.270 ;
        RECT 125.470 -12.320 125.920 -12.220 ;
        RECT 132.210 -12.220 133.360 -12.140 ;
        RECT 138.270 -11.840 139.420 -11.760 ;
        RECT 145.710 -11.760 146.160 -11.660 ;
        RECT 152.470 -8.710 152.920 -8.610 ;
        RECT 159.210 -8.610 160.360 -8.530 ;
        RECT 165.270 -8.230 166.420 -8.150 ;
        RECT 172.710 -8.150 173.160 -8.050 ;
        RECT 179.470 -5.100 179.920 -5.000 ;
        RECT 186.210 -5.000 187.360 -4.920 ;
        RECT 192.270 -4.620 193.420 -4.540 ;
        RECT 199.710 -4.540 200.160 -4.440 ;
        RECT 206.470 -1.490 206.920 -1.390 ;
        RECT 213.210 -1.390 214.360 -1.310 ;
        RECT 213.210 -1.490 213.660 -1.390 ;
        RECT 206.470 -2.640 206.910 -1.490 ;
        RECT 213.220 -2.640 213.660 -1.490 ;
        RECT 206.470 -3.290 207.620 -2.640 ;
        RECT 212.510 -3.290 213.660 -2.640 ;
        RECT 206.470 -4.440 206.910 -3.290 ;
        RECT 213.220 -4.440 213.660 -3.290 ;
        RECT 206.470 -4.540 206.920 -4.440 ;
        RECT 193.670 -4.620 194.080 -4.560 ;
        RECT 192.270 -4.920 194.080 -4.620 ;
        RECT 192.270 -5.000 193.420 -4.920 ;
        RECT 193.670 -4.980 194.080 -4.920 ;
        RECT 199.050 -4.620 199.460 -4.560 ;
        RECT 199.710 -4.620 200.860 -4.540 ;
        RECT 199.050 -4.920 200.860 -4.620 ;
        RECT 199.050 -4.980 199.460 -4.920 ;
        RECT 186.210 -5.100 186.660 -5.000 ;
        RECT 179.470 -6.250 179.910 -5.100 ;
        RECT 186.220 -6.250 186.660 -5.100 ;
        RECT 179.470 -6.900 180.620 -6.250 ;
        RECT 185.510 -6.900 186.660 -6.250 ;
        RECT 179.470 -8.050 179.910 -6.900 ;
        RECT 186.220 -8.050 186.660 -6.900 ;
        RECT 179.470 -8.150 179.920 -8.050 ;
        RECT 166.670 -8.230 167.080 -8.170 ;
        RECT 165.270 -8.530 167.080 -8.230 ;
        RECT 165.270 -8.610 166.420 -8.530 ;
        RECT 166.670 -8.590 167.080 -8.530 ;
        RECT 172.050 -8.230 172.460 -8.170 ;
        RECT 172.710 -8.230 173.860 -8.150 ;
        RECT 172.050 -8.530 173.860 -8.230 ;
        RECT 172.050 -8.590 172.460 -8.530 ;
        RECT 159.210 -8.710 159.660 -8.610 ;
        RECT 152.470 -9.860 152.910 -8.710 ;
        RECT 159.220 -9.860 159.660 -8.710 ;
        RECT 152.470 -10.510 153.620 -9.860 ;
        RECT 158.510 -10.510 159.660 -9.860 ;
        RECT 152.470 -11.660 152.910 -10.510 ;
        RECT 159.220 -11.660 159.660 -10.510 ;
        RECT 152.470 -11.760 152.920 -11.660 ;
        RECT 139.670 -11.840 140.080 -11.780 ;
        RECT 138.270 -12.140 140.080 -11.840 ;
        RECT 138.270 -12.220 139.420 -12.140 ;
        RECT 139.670 -12.200 140.080 -12.140 ;
        RECT 145.050 -11.840 145.460 -11.780 ;
        RECT 145.710 -11.840 146.860 -11.760 ;
        RECT 145.050 -12.140 146.860 -11.840 ;
        RECT 145.050 -12.200 145.460 -12.140 ;
        RECT 132.210 -12.320 132.660 -12.220 ;
        RECT 125.470 -13.470 125.910 -12.320 ;
        RECT 132.220 -13.470 132.660 -12.320 ;
        RECT 125.470 -14.120 126.620 -13.470 ;
        RECT 131.510 -14.120 132.660 -13.470 ;
        RECT 125.470 -15.270 125.910 -14.120 ;
        RECT 132.220 -15.270 132.660 -14.120 ;
        RECT 125.470 -15.370 125.920 -15.270 ;
        RECT 112.670 -15.450 113.080 -15.390 ;
        RECT 111.270 -15.750 113.080 -15.450 ;
        RECT 111.270 -15.830 112.420 -15.750 ;
        RECT 112.670 -15.810 113.080 -15.750 ;
        RECT 118.050 -15.450 118.460 -15.390 ;
        RECT 118.710 -15.450 119.860 -15.370 ;
        RECT 118.050 -15.750 119.860 -15.450 ;
        RECT 118.050 -15.810 118.460 -15.750 ;
        RECT 105.210 -15.930 105.660 -15.830 ;
        RECT 98.470 -17.080 98.910 -15.930 ;
        RECT 105.220 -17.080 105.660 -15.930 ;
        RECT 98.470 -17.730 99.620 -17.080 ;
        RECT 104.510 -17.730 105.660 -17.080 ;
        RECT 98.470 -18.880 98.910 -17.730 ;
        RECT 105.220 -18.880 105.660 -17.730 ;
        RECT 98.470 -18.980 98.920 -18.880 ;
        RECT 85.670 -19.060 86.080 -19.000 ;
        RECT 84.270 -19.360 86.080 -19.060 ;
        RECT 84.270 -19.440 85.420 -19.360 ;
        RECT 85.670 -19.420 86.080 -19.360 ;
        RECT 91.050 -19.060 91.460 -19.000 ;
        RECT 91.710 -19.060 92.860 -18.980 ;
        RECT 91.050 -19.360 92.860 -19.060 ;
        RECT 91.050 -19.420 91.460 -19.360 ;
        RECT 78.210 -19.540 78.660 -19.440 ;
        RECT 71.470 -20.690 71.910 -19.540 ;
        RECT 78.220 -20.690 78.660 -19.540 ;
        RECT 71.470 -21.340 72.620 -20.690 ;
        RECT 77.510 -21.340 78.660 -20.690 ;
        RECT 71.470 -22.490 71.910 -21.340 ;
        RECT 78.220 -22.490 78.660 -21.340 ;
        RECT 71.470 -22.590 71.920 -22.490 ;
        RECT 58.670 -22.670 59.080 -22.610 ;
        RECT 57.270 -22.970 59.080 -22.670 ;
        RECT 57.270 -23.050 58.420 -22.970 ;
        RECT 58.670 -23.030 59.080 -22.970 ;
        RECT 64.050 -22.670 64.460 -22.610 ;
        RECT 64.710 -22.670 65.860 -22.590 ;
        RECT 64.050 -22.970 65.860 -22.670 ;
        RECT 64.050 -23.030 64.460 -22.970 ;
        RECT 51.210 -23.150 51.660 -23.050 ;
        RECT 44.470 -24.300 44.910 -23.150 ;
        RECT 51.220 -24.300 51.660 -23.150 ;
        RECT 44.470 -24.950 45.620 -24.300 ;
        RECT 50.510 -24.950 51.660 -24.300 ;
        RECT 44.470 -26.100 44.910 -24.950 ;
        RECT 51.220 -26.100 51.660 -24.950 ;
        RECT 44.470 -26.200 44.920 -26.100 ;
        RECT 31.670 -26.280 32.080 -26.220 ;
        RECT 30.270 -26.580 32.080 -26.280 ;
        RECT 30.270 -26.660 31.420 -26.580 ;
        RECT 31.670 -26.640 32.080 -26.580 ;
        RECT 37.050 -26.280 37.460 -26.220 ;
        RECT 37.710 -26.280 38.860 -26.200 ;
        RECT 37.050 -26.580 38.860 -26.280 ;
        RECT 37.050 -26.640 37.460 -26.580 ;
        RECT 24.210 -26.760 24.660 -26.660 ;
        RECT 17.470 -27.910 17.910 -26.760 ;
        RECT 24.220 -27.910 24.660 -26.760 ;
        RECT 17.470 -28.560 18.620 -27.910 ;
        RECT 23.510 -28.560 24.660 -27.910 ;
        RECT 17.470 -29.710 17.910 -28.560 ;
        RECT 24.220 -29.710 24.660 -28.560 ;
        RECT 17.470 -29.810 17.920 -29.710 ;
        RECT 4.670 -29.890 5.080 -29.830 ;
        RECT 3.270 -30.190 5.080 -29.890 ;
        RECT 3.270 -30.270 4.420 -30.190 ;
        RECT 4.670 -30.250 5.080 -30.190 ;
        RECT 10.050 -29.890 10.460 -29.830 ;
        RECT 10.710 -29.890 11.860 -29.810 ;
        RECT 10.050 -30.190 11.860 -29.890 ;
        RECT 10.050 -30.250 10.460 -30.190 ;
        RECT 3.970 -30.370 4.420 -30.270 ;
        RECT 10.710 -30.270 11.860 -30.190 ;
        RECT 16.770 -29.890 17.920 -29.810 ;
        RECT 24.210 -29.810 24.660 -29.710 ;
        RECT 30.970 -26.760 31.420 -26.660 ;
        RECT 37.710 -26.660 38.860 -26.580 ;
        RECT 43.770 -26.280 44.920 -26.200 ;
        RECT 51.210 -26.200 51.660 -26.100 ;
        RECT 57.970 -23.150 58.420 -23.050 ;
        RECT 64.710 -23.050 65.860 -22.970 ;
        RECT 70.770 -22.670 71.920 -22.590 ;
        RECT 78.210 -22.590 78.660 -22.490 ;
        RECT 84.970 -19.540 85.420 -19.440 ;
        RECT 91.710 -19.440 92.860 -19.360 ;
        RECT 97.770 -19.060 98.920 -18.980 ;
        RECT 105.210 -18.980 105.660 -18.880 ;
        RECT 111.970 -15.930 112.420 -15.830 ;
        RECT 118.710 -15.830 119.860 -15.750 ;
        RECT 124.770 -15.450 125.920 -15.370 ;
        RECT 132.210 -15.370 132.660 -15.270 ;
        RECT 138.970 -12.320 139.420 -12.220 ;
        RECT 145.710 -12.220 146.860 -12.140 ;
        RECT 151.770 -11.840 152.920 -11.760 ;
        RECT 159.210 -11.760 159.660 -11.660 ;
        RECT 165.970 -8.710 166.420 -8.610 ;
        RECT 172.710 -8.610 173.860 -8.530 ;
        RECT 178.770 -8.230 179.920 -8.150 ;
        RECT 186.210 -8.150 186.660 -8.050 ;
        RECT 192.970 -5.100 193.420 -5.000 ;
        RECT 199.710 -5.000 200.860 -4.920 ;
        RECT 205.770 -4.620 206.920 -4.540 ;
        RECT 213.210 -4.540 213.660 -4.440 ;
        RECT 207.170 -4.620 207.580 -4.560 ;
        RECT 205.770 -4.920 207.580 -4.620 ;
        RECT 205.770 -5.000 206.920 -4.920 ;
        RECT 207.170 -4.980 207.580 -4.920 ;
        RECT 212.550 -4.620 212.960 -4.560 ;
        RECT 213.210 -4.620 214.360 -4.540 ;
        RECT 212.550 -4.920 214.360 -4.620 ;
        RECT 212.550 -4.980 212.960 -4.920 ;
        RECT 199.710 -5.100 200.160 -5.000 ;
        RECT 192.970 -6.250 193.410 -5.100 ;
        RECT 199.720 -6.250 200.160 -5.100 ;
        RECT 192.970 -6.900 194.120 -6.250 ;
        RECT 199.010 -6.900 200.160 -6.250 ;
        RECT 192.970 -8.050 193.410 -6.900 ;
        RECT 199.720 -8.050 200.160 -6.900 ;
        RECT 192.970 -8.150 193.420 -8.050 ;
        RECT 180.170 -8.230 180.580 -8.170 ;
        RECT 178.770 -8.530 180.580 -8.230 ;
        RECT 178.770 -8.610 179.920 -8.530 ;
        RECT 180.170 -8.590 180.580 -8.530 ;
        RECT 185.550 -8.230 185.960 -8.170 ;
        RECT 186.210 -8.230 187.360 -8.150 ;
        RECT 185.550 -8.530 187.360 -8.230 ;
        RECT 185.550 -8.590 185.960 -8.530 ;
        RECT 172.710 -8.710 173.160 -8.610 ;
        RECT 165.970 -9.860 166.410 -8.710 ;
        RECT 172.720 -9.860 173.160 -8.710 ;
        RECT 165.970 -10.510 167.120 -9.860 ;
        RECT 172.010 -10.510 173.160 -9.860 ;
        RECT 165.970 -11.660 166.410 -10.510 ;
        RECT 172.720 -11.660 173.160 -10.510 ;
        RECT 165.970 -11.760 166.420 -11.660 ;
        RECT 153.170 -11.840 153.580 -11.780 ;
        RECT 151.770 -12.140 153.580 -11.840 ;
        RECT 151.770 -12.220 152.920 -12.140 ;
        RECT 153.170 -12.200 153.580 -12.140 ;
        RECT 158.550 -11.840 158.960 -11.780 ;
        RECT 159.210 -11.840 160.360 -11.760 ;
        RECT 158.550 -12.140 160.360 -11.840 ;
        RECT 158.550 -12.200 158.960 -12.140 ;
        RECT 145.710 -12.320 146.160 -12.220 ;
        RECT 138.970 -13.470 139.410 -12.320 ;
        RECT 145.720 -13.470 146.160 -12.320 ;
        RECT 138.970 -14.120 140.120 -13.470 ;
        RECT 145.010 -14.120 146.160 -13.470 ;
        RECT 138.970 -15.270 139.410 -14.120 ;
        RECT 145.720 -15.270 146.160 -14.120 ;
        RECT 138.970 -15.370 139.420 -15.270 ;
        RECT 126.170 -15.450 126.580 -15.390 ;
        RECT 124.770 -15.750 126.580 -15.450 ;
        RECT 124.770 -15.830 125.920 -15.750 ;
        RECT 126.170 -15.810 126.580 -15.750 ;
        RECT 131.550 -15.450 131.960 -15.390 ;
        RECT 132.210 -15.450 133.360 -15.370 ;
        RECT 131.550 -15.750 133.360 -15.450 ;
        RECT 131.550 -15.810 131.960 -15.750 ;
        RECT 118.710 -15.930 119.160 -15.830 ;
        RECT 111.970 -17.080 112.410 -15.930 ;
        RECT 118.720 -17.080 119.160 -15.930 ;
        RECT 111.970 -17.730 113.120 -17.080 ;
        RECT 118.010 -17.730 119.160 -17.080 ;
        RECT 111.970 -18.880 112.410 -17.730 ;
        RECT 118.720 -18.880 119.160 -17.730 ;
        RECT 111.970 -18.980 112.420 -18.880 ;
        RECT 99.170 -19.060 99.580 -19.000 ;
        RECT 97.770 -19.360 99.580 -19.060 ;
        RECT 97.770 -19.440 98.920 -19.360 ;
        RECT 99.170 -19.420 99.580 -19.360 ;
        RECT 104.550 -19.060 104.960 -19.000 ;
        RECT 105.210 -19.060 106.360 -18.980 ;
        RECT 104.550 -19.360 106.360 -19.060 ;
        RECT 104.550 -19.420 104.960 -19.360 ;
        RECT 91.710 -19.540 92.160 -19.440 ;
        RECT 84.970 -20.690 85.410 -19.540 ;
        RECT 91.720 -20.690 92.160 -19.540 ;
        RECT 84.970 -21.340 86.120 -20.690 ;
        RECT 91.010 -21.340 92.160 -20.690 ;
        RECT 84.970 -22.490 85.410 -21.340 ;
        RECT 91.720 -22.490 92.160 -21.340 ;
        RECT 84.970 -22.590 85.420 -22.490 ;
        RECT 72.170 -22.670 72.580 -22.610 ;
        RECT 70.770 -22.970 72.580 -22.670 ;
        RECT 70.770 -23.050 71.920 -22.970 ;
        RECT 72.170 -23.030 72.580 -22.970 ;
        RECT 77.550 -22.670 77.960 -22.610 ;
        RECT 78.210 -22.670 79.360 -22.590 ;
        RECT 77.550 -22.970 79.360 -22.670 ;
        RECT 77.550 -23.030 77.960 -22.970 ;
        RECT 64.710 -23.150 65.160 -23.050 ;
        RECT 57.970 -24.300 58.410 -23.150 ;
        RECT 64.720 -24.300 65.160 -23.150 ;
        RECT 57.970 -24.950 59.120 -24.300 ;
        RECT 64.010 -24.950 65.160 -24.300 ;
        RECT 57.970 -26.100 58.410 -24.950 ;
        RECT 64.720 -26.100 65.160 -24.950 ;
        RECT 57.970 -26.200 58.420 -26.100 ;
        RECT 45.170 -26.280 45.580 -26.220 ;
        RECT 43.770 -26.580 45.580 -26.280 ;
        RECT 43.770 -26.660 44.920 -26.580 ;
        RECT 45.170 -26.640 45.580 -26.580 ;
        RECT 50.550 -26.280 50.960 -26.220 ;
        RECT 51.210 -26.280 52.360 -26.200 ;
        RECT 50.550 -26.580 52.360 -26.280 ;
        RECT 50.550 -26.640 50.960 -26.580 ;
        RECT 37.710 -26.760 38.160 -26.660 ;
        RECT 30.970 -27.910 31.410 -26.760 ;
        RECT 37.720 -27.910 38.160 -26.760 ;
        RECT 30.970 -28.560 32.120 -27.910 ;
        RECT 37.010 -28.560 38.160 -27.910 ;
        RECT 30.970 -29.710 31.410 -28.560 ;
        RECT 37.720 -29.710 38.160 -28.560 ;
        RECT 30.970 -29.810 31.420 -29.710 ;
        RECT 18.170 -29.890 18.580 -29.830 ;
        RECT 16.770 -30.190 18.580 -29.890 ;
        RECT 16.770 -30.270 17.920 -30.190 ;
        RECT 18.170 -30.250 18.580 -30.190 ;
        RECT 23.550 -29.890 23.960 -29.830 ;
        RECT 24.210 -29.890 25.360 -29.810 ;
        RECT 23.550 -30.190 25.360 -29.890 ;
        RECT 23.550 -30.250 23.960 -30.190 ;
        RECT 10.710 -30.370 11.160 -30.270 ;
        RECT 3.970 -31.520 4.410 -30.370 ;
        RECT 10.720 -31.520 11.160 -30.370 ;
        RECT 3.970 -32.170 5.120 -31.520 ;
        RECT 10.010 -32.170 11.160 -31.520 ;
        RECT 3.970 -33.320 4.410 -32.170 ;
        RECT 10.720 -33.320 11.160 -32.170 ;
        RECT 3.970 -33.420 4.420 -33.320 ;
        RECT 3.270 -33.500 4.420 -33.420 ;
        RECT 10.710 -33.420 11.160 -33.320 ;
        RECT 17.470 -30.370 17.920 -30.270 ;
        RECT 24.210 -30.270 25.360 -30.190 ;
        RECT 30.270 -29.890 31.420 -29.810 ;
        RECT 37.710 -29.810 38.160 -29.710 ;
        RECT 44.470 -26.760 44.920 -26.660 ;
        RECT 51.210 -26.660 52.360 -26.580 ;
        RECT 57.270 -26.280 58.420 -26.200 ;
        RECT 64.710 -26.200 65.160 -26.100 ;
        RECT 71.470 -23.150 71.920 -23.050 ;
        RECT 78.210 -23.050 79.360 -22.970 ;
        RECT 84.270 -22.670 85.420 -22.590 ;
        RECT 91.710 -22.590 92.160 -22.490 ;
        RECT 98.470 -19.540 98.920 -19.440 ;
        RECT 105.210 -19.440 106.360 -19.360 ;
        RECT 111.270 -19.060 112.420 -18.980 ;
        RECT 118.710 -18.980 119.160 -18.880 ;
        RECT 125.470 -15.930 125.920 -15.830 ;
        RECT 132.210 -15.830 133.360 -15.750 ;
        RECT 138.270 -15.450 139.420 -15.370 ;
        RECT 145.710 -15.370 146.160 -15.270 ;
        RECT 152.470 -12.320 152.920 -12.220 ;
        RECT 159.210 -12.220 160.360 -12.140 ;
        RECT 165.270 -11.840 166.420 -11.760 ;
        RECT 172.710 -11.760 173.160 -11.660 ;
        RECT 179.470 -8.710 179.920 -8.610 ;
        RECT 186.210 -8.610 187.360 -8.530 ;
        RECT 192.270 -8.230 193.420 -8.150 ;
        RECT 199.710 -8.150 200.160 -8.050 ;
        RECT 206.470 -5.100 206.920 -5.000 ;
        RECT 213.210 -5.000 214.360 -4.920 ;
        RECT 213.210 -5.100 213.660 -5.000 ;
        RECT 206.470 -6.250 206.910 -5.100 ;
        RECT 213.220 -6.250 213.660 -5.100 ;
        RECT 206.470 -6.900 207.620 -6.250 ;
        RECT 212.510 -6.900 213.660 -6.250 ;
        RECT 206.470 -8.050 206.910 -6.900 ;
        RECT 213.220 -8.050 213.660 -6.900 ;
        RECT 206.470 -8.150 206.920 -8.050 ;
        RECT 193.670 -8.230 194.080 -8.170 ;
        RECT 192.270 -8.530 194.080 -8.230 ;
        RECT 192.270 -8.610 193.420 -8.530 ;
        RECT 193.670 -8.590 194.080 -8.530 ;
        RECT 199.050 -8.230 199.460 -8.170 ;
        RECT 199.710 -8.230 200.860 -8.150 ;
        RECT 199.050 -8.530 200.860 -8.230 ;
        RECT 199.050 -8.590 199.460 -8.530 ;
        RECT 186.210 -8.710 186.660 -8.610 ;
        RECT 179.470 -9.860 179.910 -8.710 ;
        RECT 186.220 -9.860 186.660 -8.710 ;
        RECT 179.470 -10.510 180.620 -9.860 ;
        RECT 185.510 -10.510 186.660 -9.860 ;
        RECT 179.470 -11.660 179.910 -10.510 ;
        RECT 186.220 -11.660 186.660 -10.510 ;
        RECT 179.470 -11.760 179.920 -11.660 ;
        RECT 166.670 -11.840 167.080 -11.780 ;
        RECT 165.270 -12.140 167.080 -11.840 ;
        RECT 165.270 -12.220 166.420 -12.140 ;
        RECT 166.670 -12.200 167.080 -12.140 ;
        RECT 172.050 -11.840 172.460 -11.780 ;
        RECT 172.710 -11.840 173.860 -11.760 ;
        RECT 172.050 -12.140 173.860 -11.840 ;
        RECT 172.050 -12.200 172.460 -12.140 ;
        RECT 159.210 -12.320 159.660 -12.220 ;
        RECT 152.470 -13.470 152.910 -12.320 ;
        RECT 159.220 -13.470 159.660 -12.320 ;
        RECT 152.470 -14.120 153.620 -13.470 ;
        RECT 158.510 -14.120 159.660 -13.470 ;
        RECT 152.470 -15.270 152.910 -14.120 ;
        RECT 159.220 -15.270 159.660 -14.120 ;
        RECT 152.470 -15.370 152.920 -15.270 ;
        RECT 139.670 -15.450 140.080 -15.390 ;
        RECT 138.270 -15.750 140.080 -15.450 ;
        RECT 138.270 -15.830 139.420 -15.750 ;
        RECT 139.670 -15.810 140.080 -15.750 ;
        RECT 145.050 -15.450 145.460 -15.390 ;
        RECT 145.710 -15.450 146.860 -15.370 ;
        RECT 145.050 -15.750 146.860 -15.450 ;
        RECT 145.050 -15.810 145.460 -15.750 ;
        RECT 132.210 -15.930 132.660 -15.830 ;
        RECT 125.470 -17.080 125.910 -15.930 ;
        RECT 132.220 -17.080 132.660 -15.930 ;
        RECT 125.470 -17.730 126.620 -17.080 ;
        RECT 131.510 -17.730 132.660 -17.080 ;
        RECT 125.470 -18.880 125.910 -17.730 ;
        RECT 132.220 -18.880 132.660 -17.730 ;
        RECT 125.470 -18.980 125.920 -18.880 ;
        RECT 112.670 -19.060 113.080 -19.000 ;
        RECT 111.270 -19.360 113.080 -19.060 ;
        RECT 111.270 -19.440 112.420 -19.360 ;
        RECT 112.670 -19.420 113.080 -19.360 ;
        RECT 118.050 -19.060 118.460 -19.000 ;
        RECT 118.710 -19.060 119.860 -18.980 ;
        RECT 118.050 -19.360 119.860 -19.060 ;
        RECT 118.050 -19.420 118.460 -19.360 ;
        RECT 105.210 -19.540 105.660 -19.440 ;
        RECT 98.470 -20.690 98.910 -19.540 ;
        RECT 105.220 -20.690 105.660 -19.540 ;
        RECT 98.470 -21.340 99.620 -20.690 ;
        RECT 104.510 -21.340 105.660 -20.690 ;
        RECT 98.470 -22.490 98.910 -21.340 ;
        RECT 105.220 -22.490 105.660 -21.340 ;
        RECT 98.470 -22.590 98.920 -22.490 ;
        RECT 85.670 -22.670 86.080 -22.610 ;
        RECT 84.270 -22.970 86.080 -22.670 ;
        RECT 84.270 -23.050 85.420 -22.970 ;
        RECT 85.670 -23.030 86.080 -22.970 ;
        RECT 91.050 -22.670 91.460 -22.610 ;
        RECT 91.710 -22.670 92.860 -22.590 ;
        RECT 91.050 -22.970 92.860 -22.670 ;
        RECT 91.050 -23.030 91.460 -22.970 ;
        RECT 78.210 -23.150 78.660 -23.050 ;
        RECT 71.470 -24.300 71.910 -23.150 ;
        RECT 78.220 -24.300 78.660 -23.150 ;
        RECT 71.470 -24.950 72.620 -24.300 ;
        RECT 77.510 -24.950 78.660 -24.300 ;
        RECT 71.470 -26.100 71.910 -24.950 ;
        RECT 78.220 -26.100 78.660 -24.950 ;
        RECT 71.470 -26.200 71.920 -26.100 ;
        RECT 58.670 -26.280 59.080 -26.220 ;
        RECT 57.270 -26.580 59.080 -26.280 ;
        RECT 57.270 -26.660 58.420 -26.580 ;
        RECT 58.670 -26.640 59.080 -26.580 ;
        RECT 64.050 -26.280 64.460 -26.220 ;
        RECT 64.710 -26.280 65.860 -26.200 ;
        RECT 64.050 -26.580 65.860 -26.280 ;
        RECT 64.050 -26.640 64.460 -26.580 ;
        RECT 51.210 -26.760 51.660 -26.660 ;
        RECT 44.470 -27.910 44.910 -26.760 ;
        RECT 51.220 -27.910 51.660 -26.760 ;
        RECT 44.470 -28.560 45.620 -27.910 ;
        RECT 50.510 -28.560 51.660 -27.910 ;
        RECT 44.470 -29.710 44.910 -28.560 ;
        RECT 51.220 -29.710 51.660 -28.560 ;
        RECT 44.470 -29.810 44.920 -29.710 ;
        RECT 31.670 -29.890 32.080 -29.830 ;
        RECT 30.270 -30.190 32.080 -29.890 ;
        RECT 30.270 -30.270 31.420 -30.190 ;
        RECT 31.670 -30.250 32.080 -30.190 ;
        RECT 37.050 -29.890 37.460 -29.830 ;
        RECT 37.710 -29.890 38.860 -29.810 ;
        RECT 37.050 -30.190 38.860 -29.890 ;
        RECT 37.050 -30.250 37.460 -30.190 ;
        RECT 24.210 -30.370 24.660 -30.270 ;
        RECT 17.470 -31.520 17.910 -30.370 ;
        RECT 24.220 -31.520 24.660 -30.370 ;
        RECT 17.470 -32.170 18.620 -31.520 ;
        RECT 23.510 -32.170 24.660 -31.520 ;
        RECT 17.470 -33.320 17.910 -32.170 ;
        RECT 24.220 -33.320 24.660 -32.170 ;
        RECT 17.470 -33.420 17.920 -33.320 ;
        RECT 4.670 -33.500 5.080 -33.440 ;
        RECT 3.270 -33.800 5.080 -33.500 ;
        RECT 3.270 -33.880 4.420 -33.800 ;
        RECT 4.670 -33.860 5.080 -33.800 ;
        RECT 10.050 -33.500 10.460 -33.440 ;
        RECT 10.710 -33.500 11.860 -33.420 ;
        RECT 10.050 -33.800 11.860 -33.500 ;
        RECT 10.050 -33.860 10.460 -33.800 ;
        RECT 3.970 -33.980 4.420 -33.880 ;
        RECT 10.710 -33.880 11.860 -33.800 ;
        RECT 16.770 -33.500 17.920 -33.420 ;
        RECT 24.210 -33.420 24.660 -33.320 ;
        RECT 30.970 -30.370 31.420 -30.270 ;
        RECT 37.710 -30.270 38.860 -30.190 ;
        RECT 43.770 -29.890 44.920 -29.810 ;
        RECT 51.210 -29.810 51.660 -29.710 ;
        RECT 57.970 -26.760 58.420 -26.660 ;
        RECT 64.710 -26.660 65.860 -26.580 ;
        RECT 70.770 -26.280 71.920 -26.200 ;
        RECT 78.210 -26.200 78.660 -26.100 ;
        RECT 84.970 -23.150 85.420 -23.050 ;
        RECT 91.710 -23.050 92.860 -22.970 ;
        RECT 97.770 -22.670 98.920 -22.590 ;
        RECT 105.210 -22.590 105.660 -22.490 ;
        RECT 111.970 -19.540 112.420 -19.440 ;
        RECT 118.710 -19.440 119.860 -19.360 ;
        RECT 124.770 -19.060 125.920 -18.980 ;
        RECT 132.210 -18.980 132.660 -18.880 ;
        RECT 138.970 -15.930 139.420 -15.830 ;
        RECT 145.710 -15.830 146.860 -15.750 ;
        RECT 151.770 -15.450 152.920 -15.370 ;
        RECT 159.210 -15.370 159.660 -15.270 ;
        RECT 165.970 -12.320 166.420 -12.220 ;
        RECT 172.710 -12.220 173.860 -12.140 ;
        RECT 178.770 -11.840 179.920 -11.760 ;
        RECT 186.210 -11.760 186.660 -11.660 ;
        RECT 192.970 -8.710 193.420 -8.610 ;
        RECT 199.710 -8.610 200.860 -8.530 ;
        RECT 205.770 -8.230 206.920 -8.150 ;
        RECT 213.210 -8.150 213.660 -8.050 ;
        RECT 207.170 -8.230 207.580 -8.170 ;
        RECT 205.770 -8.530 207.580 -8.230 ;
        RECT 205.770 -8.610 206.920 -8.530 ;
        RECT 207.170 -8.590 207.580 -8.530 ;
        RECT 212.550 -8.230 212.960 -8.170 ;
        RECT 213.210 -8.230 214.360 -8.150 ;
        RECT 212.550 -8.530 214.360 -8.230 ;
        RECT 212.550 -8.590 212.960 -8.530 ;
        RECT 199.710 -8.710 200.160 -8.610 ;
        RECT 192.970 -9.860 193.410 -8.710 ;
        RECT 199.720 -9.860 200.160 -8.710 ;
        RECT 192.970 -10.510 194.120 -9.860 ;
        RECT 199.010 -10.510 200.160 -9.860 ;
        RECT 192.970 -11.660 193.410 -10.510 ;
        RECT 199.720 -11.660 200.160 -10.510 ;
        RECT 192.970 -11.760 193.420 -11.660 ;
        RECT 180.170 -11.840 180.580 -11.780 ;
        RECT 178.770 -12.140 180.580 -11.840 ;
        RECT 178.770 -12.220 179.920 -12.140 ;
        RECT 180.170 -12.200 180.580 -12.140 ;
        RECT 185.550 -11.840 185.960 -11.780 ;
        RECT 186.210 -11.840 187.360 -11.760 ;
        RECT 185.550 -12.140 187.360 -11.840 ;
        RECT 185.550 -12.200 185.960 -12.140 ;
        RECT 172.710 -12.320 173.160 -12.220 ;
        RECT 165.970 -13.470 166.410 -12.320 ;
        RECT 172.720 -13.470 173.160 -12.320 ;
        RECT 165.970 -14.120 167.120 -13.470 ;
        RECT 172.010 -14.120 173.160 -13.470 ;
        RECT 165.970 -15.270 166.410 -14.120 ;
        RECT 172.720 -15.270 173.160 -14.120 ;
        RECT 165.970 -15.370 166.420 -15.270 ;
        RECT 153.170 -15.450 153.580 -15.390 ;
        RECT 151.770 -15.750 153.580 -15.450 ;
        RECT 151.770 -15.830 152.920 -15.750 ;
        RECT 153.170 -15.810 153.580 -15.750 ;
        RECT 158.550 -15.450 158.960 -15.390 ;
        RECT 159.210 -15.450 160.360 -15.370 ;
        RECT 158.550 -15.750 160.360 -15.450 ;
        RECT 158.550 -15.810 158.960 -15.750 ;
        RECT 145.710 -15.930 146.160 -15.830 ;
        RECT 138.970 -17.080 139.410 -15.930 ;
        RECT 145.720 -17.080 146.160 -15.930 ;
        RECT 138.970 -17.730 140.120 -17.080 ;
        RECT 145.010 -17.730 146.160 -17.080 ;
        RECT 138.970 -18.880 139.410 -17.730 ;
        RECT 145.720 -18.880 146.160 -17.730 ;
        RECT 138.970 -18.980 139.420 -18.880 ;
        RECT 126.170 -19.060 126.580 -19.000 ;
        RECT 124.770 -19.360 126.580 -19.060 ;
        RECT 124.770 -19.440 125.920 -19.360 ;
        RECT 126.170 -19.420 126.580 -19.360 ;
        RECT 131.550 -19.060 131.960 -19.000 ;
        RECT 132.210 -19.060 133.360 -18.980 ;
        RECT 131.550 -19.360 133.360 -19.060 ;
        RECT 131.550 -19.420 131.960 -19.360 ;
        RECT 118.710 -19.540 119.160 -19.440 ;
        RECT 111.970 -20.690 112.410 -19.540 ;
        RECT 118.720 -20.690 119.160 -19.540 ;
        RECT 111.970 -21.340 113.120 -20.690 ;
        RECT 118.010 -21.340 119.160 -20.690 ;
        RECT 111.970 -22.490 112.410 -21.340 ;
        RECT 118.720 -22.490 119.160 -21.340 ;
        RECT 111.970 -22.590 112.420 -22.490 ;
        RECT 99.170 -22.670 99.580 -22.610 ;
        RECT 97.770 -22.970 99.580 -22.670 ;
        RECT 97.770 -23.050 98.920 -22.970 ;
        RECT 99.170 -23.030 99.580 -22.970 ;
        RECT 104.550 -22.670 104.960 -22.610 ;
        RECT 105.210 -22.670 106.360 -22.590 ;
        RECT 104.550 -22.970 106.360 -22.670 ;
        RECT 104.550 -23.030 104.960 -22.970 ;
        RECT 91.710 -23.150 92.160 -23.050 ;
        RECT 84.970 -24.300 85.410 -23.150 ;
        RECT 91.720 -24.300 92.160 -23.150 ;
        RECT 84.970 -24.950 86.120 -24.300 ;
        RECT 91.010 -24.950 92.160 -24.300 ;
        RECT 84.970 -26.100 85.410 -24.950 ;
        RECT 91.720 -26.100 92.160 -24.950 ;
        RECT 84.970 -26.200 85.420 -26.100 ;
        RECT 72.170 -26.280 72.580 -26.220 ;
        RECT 70.770 -26.580 72.580 -26.280 ;
        RECT 70.770 -26.660 71.920 -26.580 ;
        RECT 72.170 -26.640 72.580 -26.580 ;
        RECT 77.550 -26.280 77.960 -26.220 ;
        RECT 78.210 -26.280 79.360 -26.200 ;
        RECT 77.550 -26.580 79.360 -26.280 ;
        RECT 77.550 -26.640 77.960 -26.580 ;
        RECT 64.710 -26.760 65.160 -26.660 ;
        RECT 57.970 -27.910 58.410 -26.760 ;
        RECT 64.720 -27.910 65.160 -26.760 ;
        RECT 57.970 -28.560 59.120 -27.910 ;
        RECT 64.010 -28.560 65.160 -27.910 ;
        RECT 57.970 -29.710 58.410 -28.560 ;
        RECT 64.720 -29.710 65.160 -28.560 ;
        RECT 57.970 -29.810 58.420 -29.710 ;
        RECT 45.170 -29.890 45.580 -29.830 ;
        RECT 43.770 -30.190 45.580 -29.890 ;
        RECT 43.770 -30.270 44.920 -30.190 ;
        RECT 45.170 -30.250 45.580 -30.190 ;
        RECT 50.550 -29.890 50.960 -29.830 ;
        RECT 51.210 -29.890 52.360 -29.810 ;
        RECT 50.550 -30.190 52.360 -29.890 ;
        RECT 50.550 -30.250 50.960 -30.190 ;
        RECT 37.710 -30.370 38.160 -30.270 ;
        RECT 30.970 -31.520 31.410 -30.370 ;
        RECT 37.720 -31.520 38.160 -30.370 ;
        RECT 30.970 -32.170 32.120 -31.520 ;
        RECT 37.010 -32.170 38.160 -31.520 ;
        RECT 30.970 -33.320 31.410 -32.170 ;
        RECT 37.720 -33.320 38.160 -32.170 ;
        RECT 30.970 -33.420 31.420 -33.320 ;
        RECT 18.170 -33.500 18.580 -33.440 ;
        RECT 16.770 -33.800 18.580 -33.500 ;
        RECT 16.770 -33.880 17.920 -33.800 ;
        RECT 18.170 -33.860 18.580 -33.800 ;
        RECT 23.550 -33.500 23.960 -33.440 ;
        RECT 24.210 -33.500 25.360 -33.420 ;
        RECT 23.550 -33.800 25.360 -33.500 ;
        RECT 23.550 -33.860 23.960 -33.800 ;
        RECT 10.710 -33.980 11.160 -33.880 ;
        RECT 3.970 -35.130 4.410 -33.980 ;
        RECT 10.720 -35.130 11.160 -33.980 ;
        RECT 3.970 -35.780 5.120 -35.130 ;
        RECT 10.010 -35.780 11.160 -35.130 ;
        RECT 3.970 -36.930 4.410 -35.780 ;
        RECT 10.720 -36.930 11.160 -35.780 ;
        RECT 3.970 -37.030 4.420 -36.930 ;
        RECT 3.270 -37.110 4.420 -37.030 ;
        RECT 10.710 -37.030 11.160 -36.930 ;
        RECT 17.470 -33.980 17.920 -33.880 ;
        RECT 24.210 -33.880 25.360 -33.800 ;
        RECT 30.270 -33.500 31.420 -33.420 ;
        RECT 37.710 -33.420 38.160 -33.320 ;
        RECT 44.470 -30.370 44.920 -30.270 ;
        RECT 51.210 -30.270 52.360 -30.190 ;
        RECT 57.270 -29.890 58.420 -29.810 ;
        RECT 64.710 -29.810 65.160 -29.710 ;
        RECT 71.470 -26.760 71.920 -26.660 ;
        RECT 78.210 -26.660 79.360 -26.580 ;
        RECT 84.270 -26.280 85.420 -26.200 ;
        RECT 91.710 -26.200 92.160 -26.100 ;
        RECT 98.470 -23.150 98.920 -23.050 ;
        RECT 105.210 -23.050 106.360 -22.970 ;
        RECT 111.270 -22.670 112.420 -22.590 ;
        RECT 118.710 -22.590 119.160 -22.490 ;
        RECT 125.470 -19.540 125.920 -19.440 ;
        RECT 132.210 -19.440 133.360 -19.360 ;
        RECT 138.270 -19.060 139.420 -18.980 ;
        RECT 145.710 -18.980 146.160 -18.880 ;
        RECT 152.470 -15.930 152.920 -15.830 ;
        RECT 159.210 -15.830 160.360 -15.750 ;
        RECT 165.270 -15.450 166.420 -15.370 ;
        RECT 172.710 -15.370 173.160 -15.270 ;
        RECT 179.470 -12.320 179.920 -12.220 ;
        RECT 186.210 -12.220 187.360 -12.140 ;
        RECT 192.270 -11.840 193.420 -11.760 ;
        RECT 199.710 -11.760 200.160 -11.660 ;
        RECT 206.470 -8.710 206.920 -8.610 ;
        RECT 213.210 -8.610 214.360 -8.530 ;
        RECT 213.210 -8.710 213.660 -8.610 ;
        RECT 206.470 -9.860 206.910 -8.710 ;
        RECT 213.220 -9.860 213.660 -8.710 ;
        RECT 206.470 -10.510 207.620 -9.860 ;
        RECT 212.510 -10.510 213.660 -9.860 ;
        RECT 206.470 -11.660 206.910 -10.510 ;
        RECT 213.220 -11.660 213.660 -10.510 ;
        RECT 206.470 -11.760 206.920 -11.660 ;
        RECT 193.670 -11.840 194.080 -11.780 ;
        RECT 192.270 -12.140 194.080 -11.840 ;
        RECT 192.270 -12.220 193.420 -12.140 ;
        RECT 193.670 -12.200 194.080 -12.140 ;
        RECT 199.050 -11.840 199.460 -11.780 ;
        RECT 199.710 -11.840 200.860 -11.760 ;
        RECT 199.050 -12.140 200.860 -11.840 ;
        RECT 199.050 -12.200 199.460 -12.140 ;
        RECT 186.210 -12.320 186.660 -12.220 ;
        RECT 179.470 -13.470 179.910 -12.320 ;
        RECT 186.220 -13.470 186.660 -12.320 ;
        RECT 179.470 -14.120 180.620 -13.470 ;
        RECT 185.510 -14.120 186.660 -13.470 ;
        RECT 179.470 -15.270 179.910 -14.120 ;
        RECT 186.220 -15.270 186.660 -14.120 ;
        RECT 179.470 -15.370 179.920 -15.270 ;
        RECT 166.670 -15.450 167.080 -15.390 ;
        RECT 165.270 -15.750 167.080 -15.450 ;
        RECT 165.270 -15.830 166.420 -15.750 ;
        RECT 166.670 -15.810 167.080 -15.750 ;
        RECT 172.050 -15.450 172.460 -15.390 ;
        RECT 172.710 -15.450 173.860 -15.370 ;
        RECT 172.050 -15.750 173.860 -15.450 ;
        RECT 172.050 -15.810 172.460 -15.750 ;
        RECT 159.210 -15.930 159.660 -15.830 ;
        RECT 152.470 -17.080 152.910 -15.930 ;
        RECT 159.220 -17.080 159.660 -15.930 ;
        RECT 152.470 -17.730 153.620 -17.080 ;
        RECT 158.510 -17.730 159.660 -17.080 ;
        RECT 152.470 -18.880 152.910 -17.730 ;
        RECT 159.220 -18.880 159.660 -17.730 ;
        RECT 152.470 -18.980 152.920 -18.880 ;
        RECT 139.670 -19.060 140.080 -19.000 ;
        RECT 138.270 -19.360 140.080 -19.060 ;
        RECT 138.270 -19.440 139.420 -19.360 ;
        RECT 139.670 -19.420 140.080 -19.360 ;
        RECT 145.050 -19.060 145.460 -19.000 ;
        RECT 145.710 -19.060 146.860 -18.980 ;
        RECT 145.050 -19.360 146.860 -19.060 ;
        RECT 145.050 -19.420 145.460 -19.360 ;
        RECT 132.210 -19.540 132.660 -19.440 ;
        RECT 125.470 -20.690 125.910 -19.540 ;
        RECT 132.220 -20.690 132.660 -19.540 ;
        RECT 125.470 -21.340 126.620 -20.690 ;
        RECT 131.510 -21.340 132.660 -20.690 ;
        RECT 125.470 -22.490 125.910 -21.340 ;
        RECT 132.220 -22.490 132.660 -21.340 ;
        RECT 125.470 -22.590 125.920 -22.490 ;
        RECT 112.670 -22.670 113.080 -22.610 ;
        RECT 111.270 -22.970 113.080 -22.670 ;
        RECT 111.270 -23.050 112.420 -22.970 ;
        RECT 112.670 -23.030 113.080 -22.970 ;
        RECT 118.050 -22.670 118.460 -22.610 ;
        RECT 118.710 -22.670 119.860 -22.590 ;
        RECT 118.050 -22.970 119.860 -22.670 ;
        RECT 118.050 -23.030 118.460 -22.970 ;
        RECT 105.210 -23.150 105.660 -23.050 ;
        RECT 98.470 -24.300 98.910 -23.150 ;
        RECT 105.220 -24.300 105.660 -23.150 ;
        RECT 98.470 -24.950 99.620 -24.300 ;
        RECT 104.510 -24.950 105.660 -24.300 ;
        RECT 98.470 -26.100 98.910 -24.950 ;
        RECT 105.220 -26.100 105.660 -24.950 ;
        RECT 98.470 -26.200 98.920 -26.100 ;
        RECT 85.670 -26.280 86.080 -26.220 ;
        RECT 84.270 -26.580 86.080 -26.280 ;
        RECT 84.270 -26.660 85.420 -26.580 ;
        RECT 85.670 -26.640 86.080 -26.580 ;
        RECT 91.050 -26.280 91.460 -26.220 ;
        RECT 91.710 -26.280 92.860 -26.200 ;
        RECT 91.050 -26.580 92.860 -26.280 ;
        RECT 91.050 -26.640 91.460 -26.580 ;
        RECT 78.210 -26.760 78.660 -26.660 ;
        RECT 71.470 -27.910 71.910 -26.760 ;
        RECT 78.220 -27.910 78.660 -26.760 ;
        RECT 71.470 -28.560 72.620 -27.910 ;
        RECT 77.510 -28.560 78.660 -27.910 ;
        RECT 71.470 -29.710 71.910 -28.560 ;
        RECT 78.220 -29.710 78.660 -28.560 ;
        RECT 71.470 -29.810 71.920 -29.710 ;
        RECT 58.670 -29.890 59.080 -29.830 ;
        RECT 57.270 -30.190 59.080 -29.890 ;
        RECT 57.270 -30.270 58.420 -30.190 ;
        RECT 58.670 -30.250 59.080 -30.190 ;
        RECT 64.050 -29.890 64.460 -29.830 ;
        RECT 64.710 -29.890 65.860 -29.810 ;
        RECT 64.050 -30.190 65.860 -29.890 ;
        RECT 64.050 -30.250 64.460 -30.190 ;
        RECT 51.210 -30.370 51.660 -30.270 ;
        RECT 44.470 -31.520 44.910 -30.370 ;
        RECT 51.220 -31.520 51.660 -30.370 ;
        RECT 44.470 -32.170 45.620 -31.520 ;
        RECT 50.510 -32.170 51.660 -31.520 ;
        RECT 44.470 -33.320 44.910 -32.170 ;
        RECT 51.220 -33.320 51.660 -32.170 ;
        RECT 44.470 -33.420 44.920 -33.320 ;
        RECT 31.670 -33.500 32.080 -33.440 ;
        RECT 30.270 -33.800 32.080 -33.500 ;
        RECT 30.270 -33.880 31.420 -33.800 ;
        RECT 31.670 -33.860 32.080 -33.800 ;
        RECT 37.050 -33.500 37.460 -33.440 ;
        RECT 37.710 -33.500 38.860 -33.420 ;
        RECT 37.050 -33.800 38.860 -33.500 ;
        RECT 37.050 -33.860 37.460 -33.800 ;
        RECT 24.210 -33.980 24.660 -33.880 ;
        RECT 17.470 -35.130 17.910 -33.980 ;
        RECT 24.220 -35.130 24.660 -33.980 ;
        RECT 17.470 -35.780 18.620 -35.130 ;
        RECT 23.510 -35.780 24.660 -35.130 ;
        RECT 17.470 -36.930 17.910 -35.780 ;
        RECT 24.220 -36.930 24.660 -35.780 ;
        RECT 17.470 -37.030 17.920 -36.930 ;
        RECT 4.670 -37.110 5.080 -37.050 ;
        RECT 3.270 -37.410 5.080 -37.110 ;
        RECT 3.270 -37.490 4.420 -37.410 ;
        RECT 4.670 -37.470 5.080 -37.410 ;
        RECT 10.050 -37.110 10.460 -37.050 ;
        RECT 10.710 -37.110 11.860 -37.030 ;
        RECT 10.050 -37.410 11.860 -37.110 ;
        RECT 10.050 -37.470 10.460 -37.410 ;
        RECT 3.970 -37.590 4.420 -37.490 ;
        RECT 10.710 -37.490 11.860 -37.410 ;
        RECT 16.770 -37.110 17.920 -37.030 ;
        RECT 24.210 -37.030 24.660 -36.930 ;
        RECT 30.970 -33.980 31.420 -33.880 ;
        RECT 37.710 -33.880 38.860 -33.800 ;
        RECT 43.770 -33.500 44.920 -33.420 ;
        RECT 51.210 -33.420 51.660 -33.320 ;
        RECT 57.970 -30.370 58.420 -30.270 ;
        RECT 64.710 -30.270 65.860 -30.190 ;
        RECT 70.770 -29.890 71.920 -29.810 ;
        RECT 78.210 -29.810 78.660 -29.710 ;
        RECT 84.970 -26.760 85.420 -26.660 ;
        RECT 91.710 -26.660 92.860 -26.580 ;
        RECT 97.770 -26.280 98.920 -26.200 ;
        RECT 105.210 -26.200 105.660 -26.100 ;
        RECT 111.970 -23.150 112.420 -23.050 ;
        RECT 118.710 -23.050 119.860 -22.970 ;
        RECT 124.770 -22.670 125.920 -22.590 ;
        RECT 132.210 -22.590 132.660 -22.490 ;
        RECT 138.970 -19.540 139.420 -19.440 ;
        RECT 145.710 -19.440 146.860 -19.360 ;
        RECT 151.770 -19.060 152.920 -18.980 ;
        RECT 159.210 -18.980 159.660 -18.880 ;
        RECT 165.970 -15.930 166.420 -15.830 ;
        RECT 172.710 -15.830 173.860 -15.750 ;
        RECT 178.770 -15.450 179.920 -15.370 ;
        RECT 186.210 -15.370 186.660 -15.270 ;
        RECT 192.970 -12.320 193.420 -12.220 ;
        RECT 199.710 -12.220 200.860 -12.140 ;
        RECT 205.770 -11.840 206.920 -11.760 ;
        RECT 213.210 -11.760 213.660 -11.660 ;
        RECT 207.170 -11.840 207.580 -11.780 ;
        RECT 205.770 -12.140 207.580 -11.840 ;
        RECT 205.770 -12.220 206.920 -12.140 ;
        RECT 207.170 -12.200 207.580 -12.140 ;
        RECT 212.550 -11.840 212.960 -11.780 ;
        RECT 213.210 -11.840 214.360 -11.760 ;
        RECT 212.550 -12.140 214.360 -11.840 ;
        RECT 212.550 -12.200 212.960 -12.140 ;
        RECT 199.710 -12.320 200.160 -12.220 ;
        RECT 192.970 -13.470 193.410 -12.320 ;
        RECT 199.720 -13.470 200.160 -12.320 ;
        RECT 192.970 -14.120 194.120 -13.470 ;
        RECT 199.010 -14.120 200.160 -13.470 ;
        RECT 192.970 -15.270 193.410 -14.120 ;
        RECT 199.720 -15.270 200.160 -14.120 ;
        RECT 192.970 -15.370 193.420 -15.270 ;
        RECT 180.170 -15.450 180.580 -15.390 ;
        RECT 178.770 -15.750 180.580 -15.450 ;
        RECT 178.770 -15.830 179.920 -15.750 ;
        RECT 180.170 -15.810 180.580 -15.750 ;
        RECT 185.550 -15.450 185.960 -15.390 ;
        RECT 186.210 -15.450 187.360 -15.370 ;
        RECT 185.550 -15.750 187.360 -15.450 ;
        RECT 185.550 -15.810 185.960 -15.750 ;
        RECT 172.710 -15.930 173.160 -15.830 ;
        RECT 165.970 -17.080 166.410 -15.930 ;
        RECT 172.720 -17.080 173.160 -15.930 ;
        RECT 165.970 -17.730 167.120 -17.080 ;
        RECT 172.010 -17.730 173.160 -17.080 ;
        RECT 165.970 -18.880 166.410 -17.730 ;
        RECT 172.720 -18.880 173.160 -17.730 ;
        RECT 165.970 -18.980 166.420 -18.880 ;
        RECT 153.170 -19.060 153.580 -19.000 ;
        RECT 151.770 -19.360 153.580 -19.060 ;
        RECT 151.770 -19.440 152.920 -19.360 ;
        RECT 153.170 -19.420 153.580 -19.360 ;
        RECT 158.550 -19.060 158.960 -19.000 ;
        RECT 159.210 -19.060 160.360 -18.980 ;
        RECT 158.550 -19.360 160.360 -19.060 ;
        RECT 158.550 -19.420 158.960 -19.360 ;
        RECT 145.710 -19.540 146.160 -19.440 ;
        RECT 138.970 -20.690 139.410 -19.540 ;
        RECT 145.720 -20.690 146.160 -19.540 ;
        RECT 138.970 -21.340 140.120 -20.690 ;
        RECT 145.010 -21.340 146.160 -20.690 ;
        RECT 138.970 -22.490 139.410 -21.340 ;
        RECT 145.720 -22.490 146.160 -21.340 ;
        RECT 138.970 -22.590 139.420 -22.490 ;
        RECT 126.170 -22.670 126.580 -22.610 ;
        RECT 124.770 -22.970 126.580 -22.670 ;
        RECT 124.770 -23.050 125.920 -22.970 ;
        RECT 126.170 -23.030 126.580 -22.970 ;
        RECT 131.550 -22.670 131.960 -22.610 ;
        RECT 132.210 -22.670 133.360 -22.590 ;
        RECT 131.550 -22.970 133.360 -22.670 ;
        RECT 131.550 -23.030 131.960 -22.970 ;
        RECT 118.710 -23.150 119.160 -23.050 ;
        RECT 111.970 -24.300 112.410 -23.150 ;
        RECT 118.720 -24.300 119.160 -23.150 ;
        RECT 111.970 -24.950 113.120 -24.300 ;
        RECT 118.010 -24.950 119.160 -24.300 ;
        RECT 111.970 -26.100 112.410 -24.950 ;
        RECT 118.720 -26.100 119.160 -24.950 ;
        RECT 111.970 -26.200 112.420 -26.100 ;
        RECT 99.170 -26.280 99.580 -26.220 ;
        RECT 97.770 -26.580 99.580 -26.280 ;
        RECT 97.770 -26.660 98.920 -26.580 ;
        RECT 99.170 -26.640 99.580 -26.580 ;
        RECT 104.550 -26.280 104.960 -26.220 ;
        RECT 105.210 -26.280 106.360 -26.200 ;
        RECT 104.550 -26.580 106.360 -26.280 ;
        RECT 104.550 -26.640 104.960 -26.580 ;
        RECT 91.710 -26.760 92.160 -26.660 ;
        RECT 84.970 -27.910 85.410 -26.760 ;
        RECT 91.720 -27.910 92.160 -26.760 ;
        RECT 84.970 -28.560 86.120 -27.910 ;
        RECT 91.010 -28.560 92.160 -27.910 ;
        RECT 84.970 -29.710 85.410 -28.560 ;
        RECT 91.720 -29.710 92.160 -28.560 ;
        RECT 84.970 -29.810 85.420 -29.710 ;
        RECT 72.170 -29.890 72.580 -29.830 ;
        RECT 70.770 -30.190 72.580 -29.890 ;
        RECT 70.770 -30.270 71.920 -30.190 ;
        RECT 72.170 -30.250 72.580 -30.190 ;
        RECT 77.550 -29.890 77.960 -29.830 ;
        RECT 78.210 -29.890 79.360 -29.810 ;
        RECT 77.550 -30.190 79.360 -29.890 ;
        RECT 77.550 -30.250 77.960 -30.190 ;
        RECT 64.710 -30.370 65.160 -30.270 ;
        RECT 57.970 -31.520 58.410 -30.370 ;
        RECT 64.720 -31.520 65.160 -30.370 ;
        RECT 57.970 -32.170 59.120 -31.520 ;
        RECT 64.010 -32.170 65.160 -31.520 ;
        RECT 57.970 -33.320 58.410 -32.170 ;
        RECT 64.720 -33.320 65.160 -32.170 ;
        RECT 57.970 -33.420 58.420 -33.320 ;
        RECT 45.170 -33.500 45.580 -33.440 ;
        RECT 43.770 -33.800 45.580 -33.500 ;
        RECT 43.770 -33.880 44.920 -33.800 ;
        RECT 45.170 -33.860 45.580 -33.800 ;
        RECT 50.550 -33.500 50.960 -33.440 ;
        RECT 51.210 -33.500 52.360 -33.420 ;
        RECT 50.550 -33.800 52.360 -33.500 ;
        RECT 50.550 -33.860 50.960 -33.800 ;
        RECT 37.710 -33.980 38.160 -33.880 ;
        RECT 30.970 -35.130 31.410 -33.980 ;
        RECT 37.720 -35.130 38.160 -33.980 ;
        RECT 30.970 -35.780 32.120 -35.130 ;
        RECT 37.010 -35.780 38.160 -35.130 ;
        RECT 30.970 -36.930 31.410 -35.780 ;
        RECT 37.720 -36.930 38.160 -35.780 ;
        RECT 30.970 -37.030 31.420 -36.930 ;
        RECT 18.170 -37.110 18.580 -37.050 ;
        RECT 16.770 -37.410 18.580 -37.110 ;
        RECT 16.770 -37.490 17.920 -37.410 ;
        RECT 18.170 -37.470 18.580 -37.410 ;
        RECT 23.550 -37.110 23.960 -37.050 ;
        RECT 24.210 -37.110 25.360 -37.030 ;
        RECT 23.550 -37.410 25.360 -37.110 ;
        RECT 23.550 -37.470 23.960 -37.410 ;
        RECT 10.710 -37.590 11.160 -37.490 ;
        RECT 3.970 -38.740 4.410 -37.590 ;
        RECT 10.720 -38.740 11.160 -37.590 ;
        RECT 3.970 -39.390 5.120 -38.740 ;
        RECT 10.010 -39.390 11.160 -38.740 ;
        RECT 3.970 -40.540 4.410 -39.390 ;
        RECT 10.720 -40.540 11.160 -39.390 ;
        RECT 3.970 -40.640 4.420 -40.540 ;
        RECT 3.270 -40.720 4.420 -40.640 ;
        RECT 10.710 -40.640 11.160 -40.540 ;
        RECT 17.470 -37.590 17.920 -37.490 ;
        RECT 24.210 -37.490 25.360 -37.410 ;
        RECT 30.270 -37.110 31.420 -37.030 ;
        RECT 37.710 -37.030 38.160 -36.930 ;
        RECT 44.470 -33.980 44.920 -33.880 ;
        RECT 51.210 -33.880 52.360 -33.800 ;
        RECT 57.270 -33.500 58.420 -33.420 ;
        RECT 64.710 -33.420 65.160 -33.320 ;
        RECT 71.470 -30.370 71.920 -30.270 ;
        RECT 78.210 -30.270 79.360 -30.190 ;
        RECT 84.270 -29.890 85.420 -29.810 ;
        RECT 91.710 -29.810 92.160 -29.710 ;
        RECT 98.470 -26.760 98.920 -26.660 ;
        RECT 105.210 -26.660 106.360 -26.580 ;
        RECT 111.270 -26.280 112.420 -26.200 ;
        RECT 118.710 -26.200 119.160 -26.100 ;
        RECT 125.470 -23.150 125.920 -23.050 ;
        RECT 132.210 -23.050 133.360 -22.970 ;
        RECT 138.270 -22.670 139.420 -22.590 ;
        RECT 145.710 -22.590 146.160 -22.490 ;
        RECT 152.470 -19.540 152.920 -19.440 ;
        RECT 159.210 -19.440 160.360 -19.360 ;
        RECT 165.270 -19.060 166.420 -18.980 ;
        RECT 172.710 -18.980 173.160 -18.880 ;
        RECT 179.470 -15.930 179.920 -15.830 ;
        RECT 186.210 -15.830 187.360 -15.750 ;
        RECT 192.270 -15.450 193.420 -15.370 ;
        RECT 199.710 -15.370 200.160 -15.270 ;
        RECT 206.470 -12.320 206.920 -12.220 ;
        RECT 213.210 -12.220 214.360 -12.140 ;
        RECT 213.210 -12.320 213.660 -12.220 ;
        RECT 206.470 -13.470 206.910 -12.320 ;
        RECT 213.220 -13.470 213.660 -12.320 ;
        RECT 206.470 -14.120 207.620 -13.470 ;
        RECT 212.510 -14.120 213.660 -13.470 ;
        RECT 206.470 -15.270 206.910 -14.120 ;
        RECT 213.220 -15.270 213.660 -14.120 ;
        RECT 206.470 -15.370 206.920 -15.270 ;
        RECT 193.670 -15.450 194.080 -15.390 ;
        RECT 192.270 -15.750 194.080 -15.450 ;
        RECT 192.270 -15.830 193.420 -15.750 ;
        RECT 193.670 -15.810 194.080 -15.750 ;
        RECT 199.050 -15.450 199.460 -15.390 ;
        RECT 199.710 -15.450 200.860 -15.370 ;
        RECT 199.050 -15.750 200.860 -15.450 ;
        RECT 199.050 -15.810 199.460 -15.750 ;
        RECT 186.210 -15.930 186.660 -15.830 ;
        RECT 179.470 -17.080 179.910 -15.930 ;
        RECT 186.220 -17.080 186.660 -15.930 ;
        RECT 179.470 -17.730 180.620 -17.080 ;
        RECT 185.510 -17.730 186.660 -17.080 ;
        RECT 179.470 -18.880 179.910 -17.730 ;
        RECT 186.220 -18.880 186.660 -17.730 ;
        RECT 179.470 -18.980 179.920 -18.880 ;
        RECT 166.670 -19.060 167.080 -19.000 ;
        RECT 165.270 -19.360 167.080 -19.060 ;
        RECT 165.270 -19.440 166.420 -19.360 ;
        RECT 166.670 -19.420 167.080 -19.360 ;
        RECT 172.050 -19.060 172.460 -19.000 ;
        RECT 172.710 -19.060 173.860 -18.980 ;
        RECT 172.050 -19.360 173.860 -19.060 ;
        RECT 172.050 -19.420 172.460 -19.360 ;
        RECT 159.210 -19.540 159.660 -19.440 ;
        RECT 152.470 -20.690 152.910 -19.540 ;
        RECT 159.220 -20.690 159.660 -19.540 ;
        RECT 152.470 -21.340 153.620 -20.690 ;
        RECT 158.510 -21.340 159.660 -20.690 ;
        RECT 152.470 -22.490 152.910 -21.340 ;
        RECT 159.220 -22.490 159.660 -21.340 ;
        RECT 152.470 -22.590 152.920 -22.490 ;
        RECT 139.670 -22.670 140.080 -22.610 ;
        RECT 138.270 -22.970 140.080 -22.670 ;
        RECT 138.270 -23.050 139.420 -22.970 ;
        RECT 139.670 -23.030 140.080 -22.970 ;
        RECT 145.050 -22.670 145.460 -22.610 ;
        RECT 145.710 -22.670 146.860 -22.590 ;
        RECT 145.050 -22.970 146.860 -22.670 ;
        RECT 145.050 -23.030 145.460 -22.970 ;
        RECT 132.210 -23.150 132.660 -23.050 ;
        RECT 125.470 -24.300 125.910 -23.150 ;
        RECT 132.220 -24.300 132.660 -23.150 ;
        RECT 125.470 -24.950 126.620 -24.300 ;
        RECT 131.510 -24.950 132.660 -24.300 ;
        RECT 125.470 -26.100 125.910 -24.950 ;
        RECT 132.220 -26.100 132.660 -24.950 ;
        RECT 125.470 -26.200 125.920 -26.100 ;
        RECT 112.670 -26.280 113.080 -26.220 ;
        RECT 111.270 -26.580 113.080 -26.280 ;
        RECT 111.270 -26.660 112.420 -26.580 ;
        RECT 112.670 -26.640 113.080 -26.580 ;
        RECT 118.050 -26.280 118.460 -26.220 ;
        RECT 118.710 -26.280 119.860 -26.200 ;
        RECT 118.050 -26.580 119.860 -26.280 ;
        RECT 118.050 -26.640 118.460 -26.580 ;
        RECT 105.210 -26.760 105.660 -26.660 ;
        RECT 98.470 -27.910 98.910 -26.760 ;
        RECT 105.220 -27.910 105.660 -26.760 ;
        RECT 98.470 -28.560 99.620 -27.910 ;
        RECT 104.510 -28.560 105.660 -27.910 ;
        RECT 98.470 -29.710 98.910 -28.560 ;
        RECT 105.220 -29.710 105.660 -28.560 ;
        RECT 98.470 -29.810 98.920 -29.710 ;
        RECT 85.670 -29.890 86.080 -29.830 ;
        RECT 84.270 -30.190 86.080 -29.890 ;
        RECT 84.270 -30.270 85.420 -30.190 ;
        RECT 85.670 -30.250 86.080 -30.190 ;
        RECT 91.050 -29.890 91.460 -29.830 ;
        RECT 91.710 -29.890 92.860 -29.810 ;
        RECT 91.050 -30.190 92.860 -29.890 ;
        RECT 91.050 -30.250 91.460 -30.190 ;
        RECT 78.210 -30.370 78.660 -30.270 ;
        RECT 71.470 -31.520 71.910 -30.370 ;
        RECT 78.220 -31.520 78.660 -30.370 ;
        RECT 71.470 -32.170 72.620 -31.520 ;
        RECT 77.510 -32.170 78.660 -31.520 ;
        RECT 71.470 -33.320 71.910 -32.170 ;
        RECT 78.220 -33.320 78.660 -32.170 ;
        RECT 71.470 -33.420 71.920 -33.320 ;
        RECT 58.670 -33.500 59.080 -33.440 ;
        RECT 57.270 -33.800 59.080 -33.500 ;
        RECT 57.270 -33.880 58.420 -33.800 ;
        RECT 58.670 -33.860 59.080 -33.800 ;
        RECT 64.050 -33.500 64.460 -33.440 ;
        RECT 64.710 -33.500 65.860 -33.420 ;
        RECT 64.050 -33.800 65.860 -33.500 ;
        RECT 64.050 -33.860 64.460 -33.800 ;
        RECT 51.210 -33.980 51.660 -33.880 ;
        RECT 44.470 -35.130 44.910 -33.980 ;
        RECT 51.220 -35.130 51.660 -33.980 ;
        RECT 44.470 -35.780 45.620 -35.130 ;
        RECT 50.510 -35.780 51.660 -35.130 ;
        RECT 44.470 -36.930 44.910 -35.780 ;
        RECT 51.220 -36.930 51.660 -35.780 ;
        RECT 44.470 -37.030 44.920 -36.930 ;
        RECT 31.670 -37.110 32.080 -37.050 ;
        RECT 30.270 -37.410 32.080 -37.110 ;
        RECT 30.270 -37.490 31.420 -37.410 ;
        RECT 31.670 -37.470 32.080 -37.410 ;
        RECT 37.050 -37.110 37.460 -37.050 ;
        RECT 37.710 -37.110 38.860 -37.030 ;
        RECT 37.050 -37.410 38.860 -37.110 ;
        RECT 37.050 -37.470 37.460 -37.410 ;
        RECT 24.210 -37.590 24.660 -37.490 ;
        RECT 17.470 -38.740 17.910 -37.590 ;
        RECT 24.220 -38.740 24.660 -37.590 ;
        RECT 17.470 -39.390 18.620 -38.740 ;
        RECT 23.510 -39.390 24.660 -38.740 ;
        RECT 17.470 -40.540 17.910 -39.390 ;
        RECT 24.220 -40.540 24.660 -39.390 ;
        RECT 17.470 -40.640 17.920 -40.540 ;
        RECT 4.670 -40.720 5.080 -40.660 ;
        RECT 3.270 -40.940 5.080 -40.720 ;
        RECT 3.270 -41.090 3.720 -40.940 ;
        RECT 3.970 -40.980 5.080 -40.940 ;
        RECT 3.970 -41.090 4.420 -40.980 ;
        RECT 4.670 -41.080 5.080 -40.980 ;
        RECT 10.050 -40.720 10.460 -40.660 ;
        RECT 10.710 -40.720 11.860 -40.640 ;
        RECT 10.050 -40.940 11.860 -40.720 ;
        RECT 10.050 -40.980 11.160 -40.940 ;
        RECT 10.050 -41.080 10.460 -40.980 ;
        RECT 10.710 -41.090 11.160 -40.980 ;
        RECT 11.410 -41.090 11.860 -40.940 ;
        RECT 16.770 -40.720 17.920 -40.640 ;
        RECT 24.210 -40.640 24.660 -40.540 ;
        RECT 30.970 -37.590 31.420 -37.490 ;
        RECT 37.710 -37.490 38.860 -37.410 ;
        RECT 43.770 -37.110 44.920 -37.030 ;
        RECT 51.210 -37.030 51.660 -36.930 ;
        RECT 57.970 -33.980 58.420 -33.880 ;
        RECT 64.710 -33.880 65.860 -33.800 ;
        RECT 70.770 -33.500 71.920 -33.420 ;
        RECT 78.210 -33.420 78.660 -33.320 ;
        RECT 84.970 -30.370 85.420 -30.270 ;
        RECT 91.710 -30.270 92.860 -30.190 ;
        RECT 97.770 -29.890 98.920 -29.810 ;
        RECT 105.210 -29.810 105.660 -29.710 ;
        RECT 111.970 -26.760 112.420 -26.660 ;
        RECT 118.710 -26.660 119.860 -26.580 ;
        RECT 124.770 -26.280 125.920 -26.200 ;
        RECT 132.210 -26.200 132.660 -26.100 ;
        RECT 138.970 -23.150 139.420 -23.050 ;
        RECT 145.710 -23.050 146.860 -22.970 ;
        RECT 151.770 -22.670 152.920 -22.590 ;
        RECT 159.210 -22.590 159.660 -22.490 ;
        RECT 165.970 -19.540 166.420 -19.440 ;
        RECT 172.710 -19.440 173.860 -19.360 ;
        RECT 178.770 -19.060 179.920 -18.980 ;
        RECT 186.210 -18.980 186.660 -18.880 ;
        RECT 192.970 -15.930 193.420 -15.830 ;
        RECT 199.710 -15.830 200.860 -15.750 ;
        RECT 205.770 -15.450 206.920 -15.370 ;
        RECT 213.210 -15.370 213.660 -15.270 ;
        RECT 207.170 -15.450 207.580 -15.390 ;
        RECT 205.770 -15.750 207.580 -15.450 ;
        RECT 205.770 -15.830 206.920 -15.750 ;
        RECT 207.170 -15.810 207.580 -15.750 ;
        RECT 212.550 -15.450 212.960 -15.390 ;
        RECT 213.210 -15.450 214.360 -15.370 ;
        RECT 212.550 -15.750 214.360 -15.450 ;
        RECT 212.550 -15.810 212.960 -15.750 ;
        RECT 199.710 -15.930 200.160 -15.830 ;
        RECT 192.970 -17.080 193.410 -15.930 ;
        RECT 199.720 -17.080 200.160 -15.930 ;
        RECT 192.970 -17.730 194.120 -17.080 ;
        RECT 199.010 -17.730 200.160 -17.080 ;
        RECT 192.970 -18.880 193.410 -17.730 ;
        RECT 199.720 -18.880 200.160 -17.730 ;
        RECT 192.970 -18.980 193.420 -18.880 ;
        RECT 180.170 -19.060 180.580 -19.000 ;
        RECT 178.770 -19.360 180.580 -19.060 ;
        RECT 178.770 -19.440 179.920 -19.360 ;
        RECT 180.170 -19.420 180.580 -19.360 ;
        RECT 185.550 -19.060 185.960 -19.000 ;
        RECT 186.210 -19.060 187.360 -18.980 ;
        RECT 185.550 -19.360 187.360 -19.060 ;
        RECT 185.550 -19.420 185.960 -19.360 ;
        RECT 172.710 -19.540 173.160 -19.440 ;
        RECT 165.970 -20.690 166.410 -19.540 ;
        RECT 172.720 -20.690 173.160 -19.540 ;
        RECT 165.970 -21.340 167.120 -20.690 ;
        RECT 172.010 -21.340 173.160 -20.690 ;
        RECT 165.970 -22.490 166.410 -21.340 ;
        RECT 172.720 -22.490 173.160 -21.340 ;
        RECT 165.970 -22.590 166.420 -22.490 ;
        RECT 153.170 -22.670 153.580 -22.610 ;
        RECT 151.770 -22.970 153.580 -22.670 ;
        RECT 151.770 -23.050 152.920 -22.970 ;
        RECT 153.170 -23.030 153.580 -22.970 ;
        RECT 158.550 -22.670 158.960 -22.610 ;
        RECT 159.210 -22.670 160.360 -22.590 ;
        RECT 158.550 -22.970 160.360 -22.670 ;
        RECT 158.550 -23.030 158.960 -22.970 ;
        RECT 145.710 -23.150 146.160 -23.050 ;
        RECT 138.970 -24.300 139.410 -23.150 ;
        RECT 145.720 -24.300 146.160 -23.150 ;
        RECT 138.970 -24.950 140.120 -24.300 ;
        RECT 145.010 -24.950 146.160 -24.300 ;
        RECT 138.970 -26.100 139.410 -24.950 ;
        RECT 145.720 -26.100 146.160 -24.950 ;
        RECT 138.970 -26.200 139.420 -26.100 ;
        RECT 126.170 -26.280 126.580 -26.220 ;
        RECT 124.770 -26.580 126.580 -26.280 ;
        RECT 124.770 -26.660 125.920 -26.580 ;
        RECT 126.170 -26.640 126.580 -26.580 ;
        RECT 131.550 -26.280 131.960 -26.220 ;
        RECT 132.210 -26.280 133.360 -26.200 ;
        RECT 131.550 -26.580 133.360 -26.280 ;
        RECT 131.550 -26.640 131.960 -26.580 ;
        RECT 118.710 -26.760 119.160 -26.660 ;
        RECT 111.970 -27.910 112.410 -26.760 ;
        RECT 118.720 -27.910 119.160 -26.760 ;
        RECT 111.970 -28.560 113.120 -27.910 ;
        RECT 118.010 -28.560 119.160 -27.910 ;
        RECT 111.970 -29.710 112.410 -28.560 ;
        RECT 118.720 -29.710 119.160 -28.560 ;
        RECT 111.970 -29.810 112.420 -29.710 ;
        RECT 99.170 -29.890 99.580 -29.830 ;
        RECT 97.770 -30.190 99.580 -29.890 ;
        RECT 97.770 -30.270 98.920 -30.190 ;
        RECT 99.170 -30.250 99.580 -30.190 ;
        RECT 104.550 -29.890 104.960 -29.830 ;
        RECT 105.210 -29.890 106.360 -29.810 ;
        RECT 104.550 -30.190 106.360 -29.890 ;
        RECT 104.550 -30.250 104.960 -30.190 ;
        RECT 91.710 -30.370 92.160 -30.270 ;
        RECT 84.970 -31.520 85.410 -30.370 ;
        RECT 91.720 -31.520 92.160 -30.370 ;
        RECT 84.970 -32.170 86.120 -31.520 ;
        RECT 91.010 -32.170 92.160 -31.520 ;
        RECT 84.970 -33.320 85.410 -32.170 ;
        RECT 91.720 -33.320 92.160 -32.170 ;
        RECT 84.970 -33.420 85.420 -33.320 ;
        RECT 72.170 -33.500 72.580 -33.440 ;
        RECT 70.770 -33.800 72.580 -33.500 ;
        RECT 70.770 -33.880 71.920 -33.800 ;
        RECT 72.170 -33.860 72.580 -33.800 ;
        RECT 77.550 -33.500 77.960 -33.440 ;
        RECT 78.210 -33.500 79.360 -33.420 ;
        RECT 77.550 -33.800 79.360 -33.500 ;
        RECT 77.550 -33.860 77.960 -33.800 ;
        RECT 64.710 -33.980 65.160 -33.880 ;
        RECT 57.970 -35.130 58.410 -33.980 ;
        RECT 64.720 -35.130 65.160 -33.980 ;
        RECT 57.970 -35.780 59.120 -35.130 ;
        RECT 64.010 -35.780 65.160 -35.130 ;
        RECT 57.970 -36.930 58.410 -35.780 ;
        RECT 64.720 -36.930 65.160 -35.780 ;
        RECT 57.970 -37.030 58.420 -36.930 ;
        RECT 45.170 -37.110 45.580 -37.050 ;
        RECT 43.770 -37.410 45.580 -37.110 ;
        RECT 43.770 -37.490 44.920 -37.410 ;
        RECT 45.170 -37.470 45.580 -37.410 ;
        RECT 50.550 -37.110 50.960 -37.050 ;
        RECT 51.210 -37.110 52.360 -37.030 ;
        RECT 50.550 -37.410 52.360 -37.110 ;
        RECT 50.550 -37.470 50.960 -37.410 ;
        RECT 37.710 -37.590 38.160 -37.490 ;
        RECT 30.970 -38.740 31.410 -37.590 ;
        RECT 37.720 -38.740 38.160 -37.590 ;
        RECT 30.970 -39.390 32.120 -38.740 ;
        RECT 37.010 -39.390 38.160 -38.740 ;
        RECT 30.970 -40.540 31.410 -39.390 ;
        RECT 37.720 -40.540 38.160 -39.390 ;
        RECT 30.970 -40.640 31.420 -40.540 ;
        RECT 18.170 -40.720 18.580 -40.660 ;
        RECT 16.770 -40.940 18.580 -40.720 ;
        RECT 16.770 -41.090 17.220 -40.940 ;
        RECT 17.470 -40.980 18.580 -40.940 ;
        RECT 17.470 -41.090 17.920 -40.980 ;
        RECT 18.170 -41.080 18.580 -40.980 ;
        RECT 23.550 -40.720 23.960 -40.660 ;
        RECT 24.210 -40.720 25.360 -40.640 ;
        RECT 23.550 -40.940 25.360 -40.720 ;
        RECT 23.550 -40.980 24.660 -40.940 ;
        RECT 23.550 -41.080 23.960 -40.980 ;
        RECT 24.210 -41.090 24.660 -40.980 ;
        RECT 24.910 -41.090 25.360 -40.940 ;
        RECT 30.270 -40.720 31.420 -40.640 ;
        RECT 37.710 -40.640 38.160 -40.540 ;
        RECT 44.470 -37.590 44.920 -37.490 ;
        RECT 51.210 -37.490 52.360 -37.410 ;
        RECT 57.270 -37.110 58.420 -37.030 ;
        RECT 64.710 -37.030 65.160 -36.930 ;
        RECT 71.470 -33.980 71.920 -33.880 ;
        RECT 78.210 -33.880 79.360 -33.800 ;
        RECT 84.270 -33.500 85.420 -33.420 ;
        RECT 91.710 -33.420 92.160 -33.320 ;
        RECT 98.470 -30.370 98.920 -30.270 ;
        RECT 105.210 -30.270 106.360 -30.190 ;
        RECT 111.270 -29.890 112.420 -29.810 ;
        RECT 118.710 -29.810 119.160 -29.710 ;
        RECT 125.470 -26.760 125.920 -26.660 ;
        RECT 132.210 -26.660 133.360 -26.580 ;
        RECT 138.270 -26.280 139.420 -26.200 ;
        RECT 145.710 -26.200 146.160 -26.100 ;
        RECT 152.470 -23.150 152.920 -23.050 ;
        RECT 159.210 -23.050 160.360 -22.970 ;
        RECT 165.270 -22.670 166.420 -22.590 ;
        RECT 172.710 -22.590 173.160 -22.490 ;
        RECT 179.470 -19.540 179.920 -19.440 ;
        RECT 186.210 -19.440 187.360 -19.360 ;
        RECT 192.270 -19.060 193.420 -18.980 ;
        RECT 199.710 -18.980 200.160 -18.880 ;
        RECT 206.470 -15.930 206.920 -15.830 ;
        RECT 213.210 -15.830 214.360 -15.750 ;
        RECT 213.210 -15.930 213.660 -15.830 ;
        RECT 206.470 -17.080 206.910 -15.930 ;
        RECT 213.220 -17.080 213.660 -15.930 ;
        RECT 206.470 -17.730 207.620 -17.080 ;
        RECT 212.510 -17.730 213.660 -17.080 ;
        RECT 206.470 -18.880 206.910 -17.730 ;
        RECT 213.220 -18.880 213.660 -17.730 ;
        RECT 206.470 -18.980 206.920 -18.880 ;
        RECT 193.670 -19.060 194.080 -19.000 ;
        RECT 192.270 -19.360 194.080 -19.060 ;
        RECT 192.270 -19.440 193.420 -19.360 ;
        RECT 193.670 -19.420 194.080 -19.360 ;
        RECT 199.050 -19.060 199.460 -19.000 ;
        RECT 199.710 -19.060 200.860 -18.980 ;
        RECT 199.050 -19.360 200.860 -19.060 ;
        RECT 199.050 -19.420 199.460 -19.360 ;
        RECT 186.210 -19.540 186.660 -19.440 ;
        RECT 179.470 -20.690 179.910 -19.540 ;
        RECT 186.220 -20.690 186.660 -19.540 ;
        RECT 179.470 -21.340 180.620 -20.690 ;
        RECT 185.510 -21.340 186.660 -20.690 ;
        RECT 179.470 -22.490 179.910 -21.340 ;
        RECT 186.220 -22.490 186.660 -21.340 ;
        RECT 179.470 -22.590 179.920 -22.490 ;
        RECT 166.670 -22.670 167.080 -22.610 ;
        RECT 165.270 -22.970 167.080 -22.670 ;
        RECT 165.270 -23.050 166.420 -22.970 ;
        RECT 166.670 -23.030 167.080 -22.970 ;
        RECT 172.050 -22.670 172.460 -22.610 ;
        RECT 172.710 -22.670 173.860 -22.590 ;
        RECT 172.050 -22.970 173.860 -22.670 ;
        RECT 172.050 -23.030 172.460 -22.970 ;
        RECT 159.210 -23.150 159.660 -23.050 ;
        RECT 152.470 -24.300 152.910 -23.150 ;
        RECT 159.220 -24.300 159.660 -23.150 ;
        RECT 152.470 -24.950 153.620 -24.300 ;
        RECT 158.510 -24.950 159.660 -24.300 ;
        RECT 152.470 -26.100 152.910 -24.950 ;
        RECT 159.220 -26.100 159.660 -24.950 ;
        RECT 152.470 -26.200 152.920 -26.100 ;
        RECT 139.670 -26.280 140.080 -26.220 ;
        RECT 138.270 -26.580 140.080 -26.280 ;
        RECT 138.270 -26.660 139.420 -26.580 ;
        RECT 139.670 -26.640 140.080 -26.580 ;
        RECT 145.050 -26.280 145.460 -26.220 ;
        RECT 145.710 -26.280 146.860 -26.200 ;
        RECT 145.050 -26.580 146.860 -26.280 ;
        RECT 145.050 -26.640 145.460 -26.580 ;
        RECT 132.210 -26.760 132.660 -26.660 ;
        RECT 125.470 -27.910 125.910 -26.760 ;
        RECT 132.220 -27.910 132.660 -26.760 ;
        RECT 125.470 -28.560 126.620 -27.910 ;
        RECT 131.510 -28.560 132.660 -27.910 ;
        RECT 125.470 -29.710 125.910 -28.560 ;
        RECT 132.220 -29.710 132.660 -28.560 ;
        RECT 125.470 -29.810 125.920 -29.710 ;
        RECT 112.670 -29.890 113.080 -29.830 ;
        RECT 111.270 -30.190 113.080 -29.890 ;
        RECT 111.270 -30.270 112.420 -30.190 ;
        RECT 112.670 -30.250 113.080 -30.190 ;
        RECT 118.050 -29.890 118.460 -29.830 ;
        RECT 118.710 -29.890 119.860 -29.810 ;
        RECT 118.050 -30.190 119.860 -29.890 ;
        RECT 118.050 -30.250 118.460 -30.190 ;
        RECT 105.210 -30.370 105.660 -30.270 ;
        RECT 98.470 -31.520 98.910 -30.370 ;
        RECT 105.220 -31.520 105.660 -30.370 ;
        RECT 98.470 -32.170 99.620 -31.520 ;
        RECT 104.510 -32.170 105.660 -31.520 ;
        RECT 98.470 -33.320 98.910 -32.170 ;
        RECT 105.220 -33.320 105.660 -32.170 ;
        RECT 98.470 -33.420 98.920 -33.320 ;
        RECT 85.670 -33.500 86.080 -33.440 ;
        RECT 84.270 -33.800 86.080 -33.500 ;
        RECT 84.270 -33.880 85.420 -33.800 ;
        RECT 85.670 -33.860 86.080 -33.800 ;
        RECT 91.050 -33.500 91.460 -33.440 ;
        RECT 91.710 -33.500 92.860 -33.420 ;
        RECT 91.050 -33.800 92.860 -33.500 ;
        RECT 91.050 -33.860 91.460 -33.800 ;
        RECT 78.210 -33.980 78.660 -33.880 ;
        RECT 71.470 -35.130 71.910 -33.980 ;
        RECT 78.220 -35.130 78.660 -33.980 ;
        RECT 71.470 -35.780 72.620 -35.130 ;
        RECT 77.510 -35.780 78.660 -35.130 ;
        RECT 71.470 -36.930 71.910 -35.780 ;
        RECT 78.220 -36.930 78.660 -35.780 ;
        RECT 71.470 -37.030 71.920 -36.930 ;
        RECT 58.670 -37.110 59.080 -37.050 ;
        RECT 57.270 -37.410 59.080 -37.110 ;
        RECT 57.270 -37.490 58.420 -37.410 ;
        RECT 58.670 -37.470 59.080 -37.410 ;
        RECT 64.050 -37.110 64.460 -37.050 ;
        RECT 64.710 -37.110 65.860 -37.030 ;
        RECT 64.050 -37.410 65.860 -37.110 ;
        RECT 64.050 -37.470 64.460 -37.410 ;
        RECT 51.210 -37.590 51.660 -37.490 ;
        RECT 44.470 -38.740 44.910 -37.590 ;
        RECT 51.220 -38.740 51.660 -37.590 ;
        RECT 44.470 -39.390 45.620 -38.740 ;
        RECT 50.510 -39.390 51.660 -38.740 ;
        RECT 44.470 -40.540 44.910 -39.390 ;
        RECT 51.220 -40.540 51.660 -39.390 ;
        RECT 44.470 -40.640 44.920 -40.540 ;
        RECT 31.670 -40.720 32.080 -40.660 ;
        RECT 30.270 -40.940 32.080 -40.720 ;
        RECT 30.270 -41.090 30.720 -40.940 ;
        RECT 30.970 -40.980 32.080 -40.940 ;
        RECT 30.970 -41.090 31.420 -40.980 ;
        RECT 31.670 -41.080 32.080 -40.980 ;
        RECT 37.050 -40.720 37.460 -40.660 ;
        RECT 37.710 -40.720 38.860 -40.640 ;
        RECT 37.050 -40.940 38.860 -40.720 ;
        RECT 37.050 -40.980 38.160 -40.940 ;
        RECT 37.050 -41.080 37.460 -40.980 ;
        RECT 37.710 -41.090 38.160 -40.980 ;
        RECT 38.410 -41.090 38.860 -40.940 ;
        RECT 43.770 -40.720 44.920 -40.640 ;
        RECT 51.210 -40.640 51.660 -40.540 ;
        RECT 57.970 -37.590 58.420 -37.490 ;
        RECT 64.710 -37.490 65.860 -37.410 ;
        RECT 70.770 -37.110 71.920 -37.030 ;
        RECT 78.210 -37.030 78.660 -36.930 ;
        RECT 84.970 -33.980 85.420 -33.880 ;
        RECT 91.710 -33.880 92.860 -33.800 ;
        RECT 97.770 -33.500 98.920 -33.420 ;
        RECT 105.210 -33.420 105.660 -33.320 ;
        RECT 111.970 -30.370 112.420 -30.270 ;
        RECT 118.710 -30.270 119.860 -30.190 ;
        RECT 124.770 -29.890 125.920 -29.810 ;
        RECT 132.210 -29.810 132.660 -29.710 ;
        RECT 138.970 -26.760 139.420 -26.660 ;
        RECT 145.710 -26.660 146.860 -26.580 ;
        RECT 151.770 -26.280 152.920 -26.200 ;
        RECT 159.210 -26.200 159.660 -26.100 ;
        RECT 165.970 -23.150 166.420 -23.050 ;
        RECT 172.710 -23.050 173.860 -22.970 ;
        RECT 178.770 -22.670 179.920 -22.590 ;
        RECT 186.210 -22.590 186.660 -22.490 ;
        RECT 192.970 -19.540 193.420 -19.440 ;
        RECT 199.710 -19.440 200.860 -19.360 ;
        RECT 205.770 -19.060 206.920 -18.980 ;
        RECT 213.210 -18.980 213.660 -18.880 ;
        RECT 207.170 -19.060 207.580 -19.000 ;
        RECT 205.770 -19.360 207.580 -19.060 ;
        RECT 205.770 -19.440 206.920 -19.360 ;
        RECT 207.170 -19.420 207.580 -19.360 ;
        RECT 212.550 -19.060 212.960 -19.000 ;
        RECT 213.210 -19.060 214.360 -18.980 ;
        RECT 212.550 -19.360 214.360 -19.060 ;
        RECT 212.550 -19.420 212.960 -19.360 ;
        RECT 199.710 -19.540 200.160 -19.440 ;
        RECT 192.970 -20.690 193.410 -19.540 ;
        RECT 199.720 -20.690 200.160 -19.540 ;
        RECT 192.970 -21.340 194.120 -20.690 ;
        RECT 199.010 -21.340 200.160 -20.690 ;
        RECT 192.970 -22.490 193.410 -21.340 ;
        RECT 199.720 -22.490 200.160 -21.340 ;
        RECT 192.970 -22.590 193.420 -22.490 ;
        RECT 180.170 -22.670 180.580 -22.610 ;
        RECT 178.770 -22.970 180.580 -22.670 ;
        RECT 178.770 -23.050 179.920 -22.970 ;
        RECT 180.170 -23.030 180.580 -22.970 ;
        RECT 185.550 -22.670 185.960 -22.610 ;
        RECT 186.210 -22.670 187.360 -22.590 ;
        RECT 185.550 -22.970 187.360 -22.670 ;
        RECT 185.550 -23.030 185.960 -22.970 ;
        RECT 172.710 -23.150 173.160 -23.050 ;
        RECT 165.970 -24.300 166.410 -23.150 ;
        RECT 172.720 -24.300 173.160 -23.150 ;
        RECT 165.970 -24.950 167.120 -24.300 ;
        RECT 172.010 -24.950 173.160 -24.300 ;
        RECT 165.970 -26.100 166.410 -24.950 ;
        RECT 172.720 -26.100 173.160 -24.950 ;
        RECT 165.970 -26.200 166.420 -26.100 ;
        RECT 153.170 -26.280 153.580 -26.220 ;
        RECT 151.770 -26.580 153.580 -26.280 ;
        RECT 151.770 -26.660 152.920 -26.580 ;
        RECT 153.170 -26.640 153.580 -26.580 ;
        RECT 158.550 -26.280 158.960 -26.220 ;
        RECT 159.210 -26.280 160.360 -26.200 ;
        RECT 158.550 -26.580 160.360 -26.280 ;
        RECT 158.550 -26.640 158.960 -26.580 ;
        RECT 145.710 -26.760 146.160 -26.660 ;
        RECT 138.970 -27.910 139.410 -26.760 ;
        RECT 145.720 -27.910 146.160 -26.760 ;
        RECT 138.970 -28.560 140.120 -27.910 ;
        RECT 145.010 -28.560 146.160 -27.910 ;
        RECT 138.970 -29.710 139.410 -28.560 ;
        RECT 145.720 -29.710 146.160 -28.560 ;
        RECT 138.970 -29.810 139.420 -29.710 ;
        RECT 126.170 -29.890 126.580 -29.830 ;
        RECT 124.770 -30.190 126.580 -29.890 ;
        RECT 124.770 -30.270 125.920 -30.190 ;
        RECT 126.170 -30.250 126.580 -30.190 ;
        RECT 131.550 -29.890 131.960 -29.830 ;
        RECT 132.210 -29.890 133.360 -29.810 ;
        RECT 131.550 -30.190 133.360 -29.890 ;
        RECT 131.550 -30.250 131.960 -30.190 ;
        RECT 118.710 -30.370 119.160 -30.270 ;
        RECT 111.970 -31.520 112.410 -30.370 ;
        RECT 118.720 -31.520 119.160 -30.370 ;
        RECT 111.970 -32.170 113.120 -31.520 ;
        RECT 118.010 -32.170 119.160 -31.520 ;
        RECT 111.970 -33.320 112.410 -32.170 ;
        RECT 118.720 -33.320 119.160 -32.170 ;
        RECT 111.970 -33.420 112.420 -33.320 ;
        RECT 99.170 -33.500 99.580 -33.440 ;
        RECT 97.770 -33.800 99.580 -33.500 ;
        RECT 97.770 -33.880 98.920 -33.800 ;
        RECT 99.170 -33.860 99.580 -33.800 ;
        RECT 104.550 -33.500 104.960 -33.440 ;
        RECT 105.210 -33.500 106.360 -33.420 ;
        RECT 104.550 -33.800 106.360 -33.500 ;
        RECT 104.550 -33.860 104.960 -33.800 ;
        RECT 91.710 -33.980 92.160 -33.880 ;
        RECT 84.970 -35.130 85.410 -33.980 ;
        RECT 91.720 -35.130 92.160 -33.980 ;
        RECT 84.970 -35.780 86.120 -35.130 ;
        RECT 91.010 -35.780 92.160 -35.130 ;
        RECT 84.970 -36.930 85.410 -35.780 ;
        RECT 91.720 -36.930 92.160 -35.780 ;
        RECT 84.970 -37.030 85.420 -36.930 ;
        RECT 72.170 -37.110 72.580 -37.050 ;
        RECT 70.770 -37.410 72.580 -37.110 ;
        RECT 70.770 -37.490 71.920 -37.410 ;
        RECT 72.170 -37.470 72.580 -37.410 ;
        RECT 77.550 -37.110 77.960 -37.050 ;
        RECT 78.210 -37.110 79.360 -37.030 ;
        RECT 77.550 -37.410 79.360 -37.110 ;
        RECT 77.550 -37.470 77.960 -37.410 ;
        RECT 64.710 -37.590 65.160 -37.490 ;
        RECT 57.970 -38.740 58.410 -37.590 ;
        RECT 64.720 -38.740 65.160 -37.590 ;
        RECT 57.970 -39.390 59.120 -38.740 ;
        RECT 64.010 -39.390 65.160 -38.740 ;
        RECT 57.970 -40.540 58.410 -39.390 ;
        RECT 64.720 -40.540 65.160 -39.390 ;
        RECT 57.970 -40.640 58.420 -40.540 ;
        RECT 45.170 -40.720 45.580 -40.660 ;
        RECT 43.770 -40.940 45.580 -40.720 ;
        RECT 43.770 -41.090 44.220 -40.940 ;
        RECT 44.470 -40.980 45.580 -40.940 ;
        RECT 44.470 -41.090 44.920 -40.980 ;
        RECT 45.170 -41.080 45.580 -40.980 ;
        RECT 50.550 -40.720 50.960 -40.660 ;
        RECT 51.210 -40.720 52.360 -40.640 ;
        RECT 50.550 -40.940 52.360 -40.720 ;
        RECT 50.550 -40.980 51.660 -40.940 ;
        RECT 50.550 -41.080 50.960 -40.980 ;
        RECT 51.210 -41.090 51.660 -40.980 ;
        RECT 51.910 -41.090 52.360 -40.940 ;
        RECT 57.270 -40.720 58.420 -40.640 ;
        RECT 64.710 -40.640 65.160 -40.540 ;
        RECT 71.470 -37.590 71.920 -37.490 ;
        RECT 78.210 -37.490 79.360 -37.410 ;
        RECT 84.270 -37.110 85.420 -37.030 ;
        RECT 91.710 -37.030 92.160 -36.930 ;
        RECT 98.470 -33.980 98.920 -33.880 ;
        RECT 105.210 -33.880 106.360 -33.800 ;
        RECT 111.270 -33.500 112.420 -33.420 ;
        RECT 118.710 -33.420 119.160 -33.320 ;
        RECT 125.470 -30.370 125.920 -30.270 ;
        RECT 132.210 -30.270 133.360 -30.190 ;
        RECT 138.270 -29.890 139.420 -29.810 ;
        RECT 145.710 -29.810 146.160 -29.710 ;
        RECT 152.470 -26.760 152.920 -26.660 ;
        RECT 159.210 -26.660 160.360 -26.580 ;
        RECT 165.270 -26.280 166.420 -26.200 ;
        RECT 172.710 -26.200 173.160 -26.100 ;
        RECT 179.470 -23.150 179.920 -23.050 ;
        RECT 186.210 -23.050 187.360 -22.970 ;
        RECT 192.270 -22.670 193.420 -22.590 ;
        RECT 199.710 -22.590 200.160 -22.490 ;
        RECT 206.470 -19.540 206.920 -19.440 ;
        RECT 213.210 -19.440 214.360 -19.360 ;
        RECT 213.210 -19.540 213.660 -19.440 ;
        RECT 206.470 -20.690 206.910 -19.540 ;
        RECT 213.220 -20.690 213.660 -19.540 ;
        RECT 206.470 -21.340 207.620 -20.690 ;
        RECT 212.510 -21.340 213.660 -20.690 ;
        RECT 206.470 -22.490 206.910 -21.340 ;
        RECT 213.220 -22.490 213.660 -21.340 ;
        RECT 206.470 -22.590 206.920 -22.490 ;
        RECT 193.670 -22.670 194.080 -22.610 ;
        RECT 192.270 -22.970 194.080 -22.670 ;
        RECT 192.270 -23.050 193.420 -22.970 ;
        RECT 193.670 -23.030 194.080 -22.970 ;
        RECT 199.050 -22.670 199.460 -22.610 ;
        RECT 199.710 -22.670 200.860 -22.590 ;
        RECT 199.050 -22.970 200.860 -22.670 ;
        RECT 199.050 -23.030 199.460 -22.970 ;
        RECT 186.210 -23.150 186.660 -23.050 ;
        RECT 179.470 -24.300 179.910 -23.150 ;
        RECT 186.220 -24.300 186.660 -23.150 ;
        RECT 179.470 -24.950 180.620 -24.300 ;
        RECT 185.510 -24.950 186.660 -24.300 ;
        RECT 179.470 -26.100 179.910 -24.950 ;
        RECT 186.220 -26.100 186.660 -24.950 ;
        RECT 179.470 -26.200 179.920 -26.100 ;
        RECT 166.670 -26.280 167.080 -26.220 ;
        RECT 165.270 -26.580 167.080 -26.280 ;
        RECT 165.270 -26.660 166.420 -26.580 ;
        RECT 166.670 -26.640 167.080 -26.580 ;
        RECT 172.050 -26.280 172.460 -26.220 ;
        RECT 172.710 -26.280 173.860 -26.200 ;
        RECT 172.050 -26.580 173.860 -26.280 ;
        RECT 172.050 -26.640 172.460 -26.580 ;
        RECT 159.210 -26.760 159.660 -26.660 ;
        RECT 152.470 -27.910 152.910 -26.760 ;
        RECT 159.220 -27.910 159.660 -26.760 ;
        RECT 152.470 -28.560 153.620 -27.910 ;
        RECT 158.510 -28.560 159.660 -27.910 ;
        RECT 152.470 -29.710 152.910 -28.560 ;
        RECT 159.220 -29.710 159.660 -28.560 ;
        RECT 152.470 -29.810 152.920 -29.710 ;
        RECT 139.670 -29.890 140.080 -29.830 ;
        RECT 138.270 -30.190 140.080 -29.890 ;
        RECT 138.270 -30.270 139.420 -30.190 ;
        RECT 139.670 -30.250 140.080 -30.190 ;
        RECT 145.050 -29.890 145.460 -29.830 ;
        RECT 145.710 -29.890 146.860 -29.810 ;
        RECT 145.050 -30.190 146.860 -29.890 ;
        RECT 145.050 -30.250 145.460 -30.190 ;
        RECT 132.210 -30.370 132.660 -30.270 ;
        RECT 125.470 -31.520 125.910 -30.370 ;
        RECT 132.220 -31.520 132.660 -30.370 ;
        RECT 125.470 -32.170 126.620 -31.520 ;
        RECT 131.510 -32.170 132.660 -31.520 ;
        RECT 125.470 -33.320 125.910 -32.170 ;
        RECT 132.220 -33.320 132.660 -32.170 ;
        RECT 125.470 -33.420 125.920 -33.320 ;
        RECT 112.670 -33.500 113.080 -33.440 ;
        RECT 111.270 -33.800 113.080 -33.500 ;
        RECT 111.270 -33.880 112.420 -33.800 ;
        RECT 112.670 -33.860 113.080 -33.800 ;
        RECT 118.050 -33.500 118.460 -33.440 ;
        RECT 118.710 -33.500 119.860 -33.420 ;
        RECT 118.050 -33.800 119.860 -33.500 ;
        RECT 118.050 -33.860 118.460 -33.800 ;
        RECT 105.210 -33.980 105.660 -33.880 ;
        RECT 98.470 -35.130 98.910 -33.980 ;
        RECT 105.220 -35.130 105.660 -33.980 ;
        RECT 98.470 -35.780 99.620 -35.130 ;
        RECT 104.510 -35.780 105.660 -35.130 ;
        RECT 98.470 -36.930 98.910 -35.780 ;
        RECT 105.220 -36.930 105.660 -35.780 ;
        RECT 98.470 -37.030 98.920 -36.930 ;
        RECT 85.670 -37.110 86.080 -37.050 ;
        RECT 84.270 -37.410 86.080 -37.110 ;
        RECT 84.270 -37.490 85.420 -37.410 ;
        RECT 85.670 -37.470 86.080 -37.410 ;
        RECT 91.050 -37.110 91.460 -37.050 ;
        RECT 91.710 -37.110 92.860 -37.030 ;
        RECT 91.050 -37.410 92.860 -37.110 ;
        RECT 91.050 -37.470 91.460 -37.410 ;
        RECT 78.210 -37.590 78.660 -37.490 ;
        RECT 71.470 -38.740 71.910 -37.590 ;
        RECT 78.220 -38.740 78.660 -37.590 ;
        RECT 71.470 -39.390 72.620 -38.740 ;
        RECT 77.510 -39.390 78.660 -38.740 ;
        RECT 71.470 -40.540 71.910 -39.390 ;
        RECT 78.220 -40.540 78.660 -39.390 ;
        RECT 71.470 -40.640 71.920 -40.540 ;
        RECT 58.670 -40.720 59.080 -40.660 ;
        RECT 57.270 -40.940 59.080 -40.720 ;
        RECT 57.270 -41.090 57.720 -40.940 ;
        RECT 57.970 -40.980 59.080 -40.940 ;
        RECT 57.970 -41.090 58.420 -40.980 ;
        RECT 58.670 -41.080 59.080 -40.980 ;
        RECT 64.050 -40.720 64.460 -40.660 ;
        RECT 64.710 -40.720 65.860 -40.640 ;
        RECT 64.050 -40.940 65.860 -40.720 ;
        RECT 64.050 -40.980 65.160 -40.940 ;
        RECT 64.050 -41.080 64.460 -40.980 ;
        RECT 64.710 -41.090 65.160 -40.980 ;
        RECT 65.410 -41.090 65.860 -40.940 ;
        RECT 70.770 -40.720 71.920 -40.640 ;
        RECT 78.210 -40.640 78.660 -40.540 ;
        RECT 84.970 -37.590 85.420 -37.490 ;
        RECT 91.710 -37.490 92.860 -37.410 ;
        RECT 97.770 -37.110 98.920 -37.030 ;
        RECT 105.210 -37.030 105.660 -36.930 ;
        RECT 111.970 -33.980 112.420 -33.880 ;
        RECT 118.710 -33.880 119.860 -33.800 ;
        RECT 124.770 -33.500 125.920 -33.420 ;
        RECT 132.210 -33.420 132.660 -33.320 ;
        RECT 138.970 -30.370 139.420 -30.270 ;
        RECT 145.710 -30.270 146.860 -30.190 ;
        RECT 151.770 -29.890 152.920 -29.810 ;
        RECT 159.210 -29.810 159.660 -29.710 ;
        RECT 165.970 -26.760 166.420 -26.660 ;
        RECT 172.710 -26.660 173.860 -26.580 ;
        RECT 178.770 -26.280 179.920 -26.200 ;
        RECT 186.210 -26.200 186.660 -26.100 ;
        RECT 192.970 -23.150 193.420 -23.050 ;
        RECT 199.710 -23.050 200.860 -22.970 ;
        RECT 205.770 -22.670 206.920 -22.590 ;
        RECT 213.210 -22.590 213.660 -22.490 ;
        RECT 207.170 -22.670 207.580 -22.610 ;
        RECT 205.770 -22.970 207.580 -22.670 ;
        RECT 205.770 -23.050 206.920 -22.970 ;
        RECT 207.170 -23.030 207.580 -22.970 ;
        RECT 212.550 -22.670 212.960 -22.610 ;
        RECT 213.210 -22.670 214.360 -22.590 ;
        RECT 212.550 -22.970 214.360 -22.670 ;
        RECT 212.550 -23.030 212.960 -22.970 ;
        RECT 199.710 -23.150 200.160 -23.050 ;
        RECT 192.970 -24.300 193.410 -23.150 ;
        RECT 199.720 -24.300 200.160 -23.150 ;
        RECT 192.970 -24.950 194.120 -24.300 ;
        RECT 199.010 -24.950 200.160 -24.300 ;
        RECT 192.970 -26.100 193.410 -24.950 ;
        RECT 199.720 -26.100 200.160 -24.950 ;
        RECT 192.970 -26.200 193.420 -26.100 ;
        RECT 180.170 -26.280 180.580 -26.220 ;
        RECT 178.770 -26.580 180.580 -26.280 ;
        RECT 178.770 -26.660 179.920 -26.580 ;
        RECT 180.170 -26.640 180.580 -26.580 ;
        RECT 185.550 -26.280 185.960 -26.220 ;
        RECT 186.210 -26.280 187.360 -26.200 ;
        RECT 185.550 -26.580 187.360 -26.280 ;
        RECT 185.550 -26.640 185.960 -26.580 ;
        RECT 172.710 -26.760 173.160 -26.660 ;
        RECT 165.970 -27.910 166.410 -26.760 ;
        RECT 172.720 -27.910 173.160 -26.760 ;
        RECT 165.970 -28.560 167.120 -27.910 ;
        RECT 172.010 -28.560 173.160 -27.910 ;
        RECT 165.970 -29.710 166.410 -28.560 ;
        RECT 172.720 -29.710 173.160 -28.560 ;
        RECT 165.970 -29.810 166.420 -29.710 ;
        RECT 153.170 -29.890 153.580 -29.830 ;
        RECT 151.770 -30.190 153.580 -29.890 ;
        RECT 151.770 -30.270 152.920 -30.190 ;
        RECT 153.170 -30.250 153.580 -30.190 ;
        RECT 158.550 -29.890 158.960 -29.830 ;
        RECT 159.210 -29.890 160.360 -29.810 ;
        RECT 158.550 -30.190 160.360 -29.890 ;
        RECT 158.550 -30.250 158.960 -30.190 ;
        RECT 145.710 -30.370 146.160 -30.270 ;
        RECT 138.970 -31.520 139.410 -30.370 ;
        RECT 145.720 -31.520 146.160 -30.370 ;
        RECT 138.970 -32.170 140.120 -31.520 ;
        RECT 145.010 -32.170 146.160 -31.520 ;
        RECT 138.970 -33.320 139.410 -32.170 ;
        RECT 145.720 -33.320 146.160 -32.170 ;
        RECT 138.970 -33.420 139.420 -33.320 ;
        RECT 126.170 -33.500 126.580 -33.440 ;
        RECT 124.770 -33.800 126.580 -33.500 ;
        RECT 124.770 -33.880 125.920 -33.800 ;
        RECT 126.170 -33.860 126.580 -33.800 ;
        RECT 131.550 -33.500 131.960 -33.440 ;
        RECT 132.210 -33.500 133.360 -33.420 ;
        RECT 131.550 -33.800 133.360 -33.500 ;
        RECT 131.550 -33.860 131.960 -33.800 ;
        RECT 118.710 -33.980 119.160 -33.880 ;
        RECT 111.970 -35.130 112.410 -33.980 ;
        RECT 118.720 -35.130 119.160 -33.980 ;
        RECT 111.970 -35.780 113.120 -35.130 ;
        RECT 118.010 -35.780 119.160 -35.130 ;
        RECT 111.970 -36.930 112.410 -35.780 ;
        RECT 118.720 -36.930 119.160 -35.780 ;
        RECT 111.970 -37.030 112.420 -36.930 ;
        RECT 99.170 -37.110 99.580 -37.050 ;
        RECT 97.770 -37.410 99.580 -37.110 ;
        RECT 97.770 -37.490 98.920 -37.410 ;
        RECT 99.170 -37.470 99.580 -37.410 ;
        RECT 104.550 -37.110 104.960 -37.050 ;
        RECT 105.210 -37.110 106.360 -37.030 ;
        RECT 104.550 -37.410 106.360 -37.110 ;
        RECT 104.550 -37.470 104.960 -37.410 ;
        RECT 91.710 -37.590 92.160 -37.490 ;
        RECT 84.970 -38.740 85.410 -37.590 ;
        RECT 91.720 -38.740 92.160 -37.590 ;
        RECT 84.970 -39.390 86.120 -38.740 ;
        RECT 91.010 -39.390 92.160 -38.740 ;
        RECT 84.970 -40.540 85.410 -39.390 ;
        RECT 91.720 -40.540 92.160 -39.390 ;
        RECT 84.970 -40.640 85.420 -40.540 ;
        RECT 72.170 -40.720 72.580 -40.660 ;
        RECT 70.770 -40.940 72.580 -40.720 ;
        RECT 70.770 -41.090 71.220 -40.940 ;
        RECT 71.470 -40.980 72.580 -40.940 ;
        RECT 71.470 -41.090 71.920 -40.980 ;
        RECT 72.170 -41.080 72.580 -40.980 ;
        RECT 77.550 -40.720 77.960 -40.660 ;
        RECT 78.210 -40.720 79.360 -40.640 ;
        RECT 77.550 -40.940 79.360 -40.720 ;
        RECT 77.550 -40.980 78.660 -40.940 ;
        RECT 77.550 -41.080 77.960 -40.980 ;
        RECT 78.210 -41.090 78.660 -40.980 ;
        RECT 78.910 -41.090 79.360 -40.940 ;
        RECT 84.270 -40.720 85.420 -40.640 ;
        RECT 91.710 -40.640 92.160 -40.540 ;
        RECT 98.470 -37.590 98.920 -37.490 ;
        RECT 105.210 -37.490 106.360 -37.410 ;
        RECT 111.270 -37.110 112.420 -37.030 ;
        RECT 118.710 -37.030 119.160 -36.930 ;
        RECT 125.470 -33.980 125.920 -33.880 ;
        RECT 132.210 -33.880 133.360 -33.800 ;
        RECT 138.270 -33.500 139.420 -33.420 ;
        RECT 145.710 -33.420 146.160 -33.320 ;
        RECT 152.470 -30.370 152.920 -30.270 ;
        RECT 159.210 -30.270 160.360 -30.190 ;
        RECT 165.270 -29.890 166.420 -29.810 ;
        RECT 172.710 -29.810 173.160 -29.710 ;
        RECT 179.470 -26.760 179.920 -26.660 ;
        RECT 186.210 -26.660 187.360 -26.580 ;
        RECT 192.270 -26.280 193.420 -26.200 ;
        RECT 199.710 -26.200 200.160 -26.100 ;
        RECT 206.470 -23.150 206.920 -23.050 ;
        RECT 213.210 -23.050 214.360 -22.970 ;
        RECT 213.210 -23.150 213.660 -23.050 ;
        RECT 206.470 -24.300 206.910 -23.150 ;
        RECT 213.220 -24.300 213.660 -23.150 ;
        RECT 206.470 -24.950 207.620 -24.300 ;
        RECT 212.510 -24.950 213.660 -24.300 ;
        RECT 206.470 -26.100 206.910 -24.950 ;
        RECT 213.220 -26.100 213.660 -24.950 ;
        RECT 206.470 -26.200 206.920 -26.100 ;
        RECT 193.670 -26.280 194.080 -26.220 ;
        RECT 192.270 -26.580 194.080 -26.280 ;
        RECT 192.270 -26.660 193.420 -26.580 ;
        RECT 193.670 -26.640 194.080 -26.580 ;
        RECT 199.050 -26.280 199.460 -26.220 ;
        RECT 199.710 -26.280 200.860 -26.200 ;
        RECT 199.050 -26.580 200.860 -26.280 ;
        RECT 199.050 -26.640 199.460 -26.580 ;
        RECT 186.210 -26.760 186.660 -26.660 ;
        RECT 179.470 -27.910 179.910 -26.760 ;
        RECT 186.220 -27.910 186.660 -26.760 ;
        RECT 179.470 -28.560 180.620 -27.910 ;
        RECT 185.510 -28.560 186.660 -27.910 ;
        RECT 179.470 -29.710 179.910 -28.560 ;
        RECT 186.220 -29.710 186.660 -28.560 ;
        RECT 179.470 -29.810 179.920 -29.710 ;
        RECT 166.670 -29.890 167.080 -29.830 ;
        RECT 165.270 -30.190 167.080 -29.890 ;
        RECT 165.270 -30.270 166.420 -30.190 ;
        RECT 166.670 -30.250 167.080 -30.190 ;
        RECT 172.050 -29.890 172.460 -29.830 ;
        RECT 172.710 -29.890 173.860 -29.810 ;
        RECT 172.050 -30.190 173.860 -29.890 ;
        RECT 172.050 -30.250 172.460 -30.190 ;
        RECT 159.210 -30.370 159.660 -30.270 ;
        RECT 152.470 -31.520 152.910 -30.370 ;
        RECT 159.220 -31.520 159.660 -30.370 ;
        RECT 152.470 -32.170 153.620 -31.520 ;
        RECT 158.510 -32.170 159.660 -31.520 ;
        RECT 152.470 -33.320 152.910 -32.170 ;
        RECT 159.220 -33.320 159.660 -32.170 ;
        RECT 152.470 -33.420 152.920 -33.320 ;
        RECT 139.670 -33.500 140.080 -33.440 ;
        RECT 138.270 -33.800 140.080 -33.500 ;
        RECT 138.270 -33.880 139.420 -33.800 ;
        RECT 139.670 -33.860 140.080 -33.800 ;
        RECT 145.050 -33.500 145.460 -33.440 ;
        RECT 145.710 -33.500 146.860 -33.420 ;
        RECT 145.050 -33.800 146.860 -33.500 ;
        RECT 145.050 -33.860 145.460 -33.800 ;
        RECT 132.210 -33.980 132.660 -33.880 ;
        RECT 125.470 -35.130 125.910 -33.980 ;
        RECT 132.220 -35.130 132.660 -33.980 ;
        RECT 125.470 -35.780 126.620 -35.130 ;
        RECT 131.510 -35.780 132.660 -35.130 ;
        RECT 125.470 -36.930 125.910 -35.780 ;
        RECT 132.220 -36.930 132.660 -35.780 ;
        RECT 125.470 -37.030 125.920 -36.930 ;
        RECT 112.670 -37.110 113.080 -37.050 ;
        RECT 111.270 -37.410 113.080 -37.110 ;
        RECT 111.270 -37.490 112.420 -37.410 ;
        RECT 112.670 -37.470 113.080 -37.410 ;
        RECT 118.050 -37.110 118.460 -37.050 ;
        RECT 118.710 -37.110 119.860 -37.030 ;
        RECT 118.050 -37.410 119.860 -37.110 ;
        RECT 118.050 -37.470 118.460 -37.410 ;
        RECT 105.210 -37.590 105.660 -37.490 ;
        RECT 98.470 -38.740 98.910 -37.590 ;
        RECT 105.220 -38.740 105.660 -37.590 ;
        RECT 98.470 -39.390 99.620 -38.740 ;
        RECT 104.510 -39.390 105.660 -38.740 ;
        RECT 98.470 -40.540 98.910 -39.390 ;
        RECT 105.220 -40.540 105.660 -39.390 ;
        RECT 98.470 -40.640 98.920 -40.540 ;
        RECT 85.670 -40.720 86.080 -40.660 ;
        RECT 84.270 -40.940 86.080 -40.720 ;
        RECT 84.270 -41.090 84.720 -40.940 ;
        RECT 84.970 -40.980 86.080 -40.940 ;
        RECT 84.970 -41.090 85.420 -40.980 ;
        RECT 85.670 -41.080 86.080 -40.980 ;
        RECT 91.050 -40.720 91.460 -40.660 ;
        RECT 91.710 -40.720 92.860 -40.640 ;
        RECT 91.050 -40.940 92.860 -40.720 ;
        RECT 91.050 -40.980 92.160 -40.940 ;
        RECT 91.050 -41.080 91.460 -40.980 ;
        RECT 91.710 -41.090 92.160 -40.980 ;
        RECT 92.410 -41.090 92.860 -40.940 ;
        RECT 97.770 -40.720 98.920 -40.640 ;
        RECT 105.210 -40.640 105.660 -40.540 ;
        RECT 111.970 -37.590 112.420 -37.490 ;
        RECT 118.710 -37.490 119.860 -37.410 ;
        RECT 124.770 -37.110 125.920 -37.030 ;
        RECT 132.210 -37.030 132.660 -36.930 ;
        RECT 138.970 -33.980 139.420 -33.880 ;
        RECT 145.710 -33.880 146.860 -33.800 ;
        RECT 151.770 -33.500 152.920 -33.420 ;
        RECT 159.210 -33.420 159.660 -33.320 ;
        RECT 165.970 -30.370 166.420 -30.270 ;
        RECT 172.710 -30.270 173.860 -30.190 ;
        RECT 178.770 -29.890 179.920 -29.810 ;
        RECT 186.210 -29.810 186.660 -29.710 ;
        RECT 192.970 -26.760 193.420 -26.660 ;
        RECT 199.710 -26.660 200.860 -26.580 ;
        RECT 205.770 -26.280 206.920 -26.200 ;
        RECT 213.210 -26.200 213.660 -26.100 ;
        RECT 207.170 -26.280 207.580 -26.220 ;
        RECT 205.770 -26.580 207.580 -26.280 ;
        RECT 205.770 -26.660 206.920 -26.580 ;
        RECT 207.170 -26.640 207.580 -26.580 ;
        RECT 212.550 -26.280 212.960 -26.220 ;
        RECT 213.210 -26.280 214.360 -26.200 ;
        RECT 212.550 -26.580 214.360 -26.280 ;
        RECT 212.550 -26.640 212.960 -26.580 ;
        RECT 199.710 -26.760 200.160 -26.660 ;
        RECT 192.970 -27.910 193.410 -26.760 ;
        RECT 199.720 -27.910 200.160 -26.760 ;
        RECT 192.970 -28.560 194.120 -27.910 ;
        RECT 199.010 -28.560 200.160 -27.910 ;
        RECT 192.970 -29.710 193.410 -28.560 ;
        RECT 199.720 -29.710 200.160 -28.560 ;
        RECT 192.970 -29.810 193.420 -29.710 ;
        RECT 180.170 -29.890 180.580 -29.830 ;
        RECT 178.770 -30.190 180.580 -29.890 ;
        RECT 178.770 -30.270 179.920 -30.190 ;
        RECT 180.170 -30.250 180.580 -30.190 ;
        RECT 185.550 -29.890 185.960 -29.830 ;
        RECT 186.210 -29.890 187.360 -29.810 ;
        RECT 185.550 -30.190 187.360 -29.890 ;
        RECT 185.550 -30.250 185.960 -30.190 ;
        RECT 172.710 -30.370 173.160 -30.270 ;
        RECT 165.970 -31.520 166.410 -30.370 ;
        RECT 172.720 -31.520 173.160 -30.370 ;
        RECT 165.970 -32.170 167.120 -31.520 ;
        RECT 172.010 -32.170 173.160 -31.520 ;
        RECT 165.970 -33.320 166.410 -32.170 ;
        RECT 172.720 -33.320 173.160 -32.170 ;
        RECT 165.970 -33.420 166.420 -33.320 ;
        RECT 153.170 -33.500 153.580 -33.440 ;
        RECT 151.770 -33.800 153.580 -33.500 ;
        RECT 151.770 -33.880 152.920 -33.800 ;
        RECT 153.170 -33.860 153.580 -33.800 ;
        RECT 158.550 -33.500 158.960 -33.440 ;
        RECT 159.210 -33.500 160.360 -33.420 ;
        RECT 158.550 -33.800 160.360 -33.500 ;
        RECT 158.550 -33.860 158.960 -33.800 ;
        RECT 145.710 -33.980 146.160 -33.880 ;
        RECT 138.970 -35.130 139.410 -33.980 ;
        RECT 145.720 -35.130 146.160 -33.980 ;
        RECT 138.970 -35.780 140.120 -35.130 ;
        RECT 145.010 -35.780 146.160 -35.130 ;
        RECT 138.970 -36.930 139.410 -35.780 ;
        RECT 145.720 -36.930 146.160 -35.780 ;
        RECT 138.970 -37.030 139.420 -36.930 ;
        RECT 126.170 -37.110 126.580 -37.050 ;
        RECT 124.770 -37.410 126.580 -37.110 ;
        RECT 124.770 -37.490 125.920 -37.410 ;
        RECT 126.170 -37.470 126.580 -37.410 ;
        RECT 131.550 -37.110 131.960 -37.050 ;
        RECT 132.210 -37.110 133.360 -37.030 ;
        RECT 131.550 -37.410 133.360 -37.110 ;
        RECT 131.550 -37.470 131.960 -37.410 ;
        RECT 118.710 -37.590 119.160 -37.490 ;
        RECT 111.970 -38.740 112.410 -37.590 ;
        RECT 118.720 -38.740 119.160 -37.590 ;
        RECT 111.970 -39.390 113.120 -38.740 ;
        RECT 118.010 -39.390 119.160 -38.740 ;
        RECT 111.970 -40.540 112.410 -39.390 ;
        RECT 118.720 -40.540 119.160 -39.390 ;
        RECT 111.970 -40.640 112.420 -40.540 ;
        RECT 99.170 -40.720 99.580 -40.660 ;
        RECT 97.770 -40.940 99.580 -40.720 ;
        RECT 97.770 -41.090 98.220 -40.940 ;
        RECT 98.470 -40.980 99.580 -40.940 ;
        RECT 98.470 -41.090 98.920 -40.980 ;
        RECT 99.170 -41.080 99.580 -40.980 ;
        RECT 104.550 -40.720 104.960 -40.660 ;
        RECT 105.210 -40.720 106.360 -40.640 ;
        RECT 104.550 -40.940 106.360 -40.720 ;
        RECT 104.550 -40.980 105.660 -40.940 ;
        RECT 104.550 -41.080 104.960 -40.980 ;
        RECT 105.210 -41.090 105.660 -40.980 ;
        RECT 105.910 -41.090 106.360 -40.940 ;
        RECT 111.270 -40.720 112.420 -40.640 ;
        RECT 118.710 -40.640 119.160 -40.540 ;
        RECT 125.470 -37.590 125.920 -37.490 ;
        RECT 132.210 -37.490 133.360 -37.410 ;
        RECT 138.270 -37.110 139.420 -37.030 ;
        RECT 145.710 -37.030 146.160 -36.930 ;
        RECT 152.470 -33.980 152.920 -33.880 ;
        RECT 159.210 -33.880 160.360 -33.800 ;
        RECT 165.270 -33.500 166.420 -33.420 ;
        RECT 172.710 -33.420 173.160 -33.320 ;
        RECT 179.470 -30.370 179.920 -30.270 ;
        RECT 186.210 -30.270 187.360 -30.190 ;
        RECT 192.270 -29.890 193.420 -29.810 ;
        RECT 199.710 -29.810 200.160 -29.710 ;
        RECT 206.470 -26.760 206.920 -26.660 ;
        RECT 213.210 -26.660 214.360 -26.580 ;
        RECT 213.210 -26.760 213.660 -26.660 ;
        RECT 206.470 -27.910 206.910 -26.760 ;
        RECT 213.220 -27.910 213.660 -26.760 ;
        RECT 206.470 -28.560 207.620 -27.910 ;
        RECT 212.510 -28.560 213.660 -27.910 ;
        RECT 206.470 -29.710 206.910 -28.560 ;
        RECT 213.220 -29.710 213.660 -28.560 ;
        RECT 206.470 -29.810 206.920 -29.710 ;
        RECT 193.670 -29.890 194.080 -29.830 ;
        RECT 192.270 -30.190 194.080 -29.890 ;
        RECT 192.270 -30.270 193.420 -30.190 ;
        RECT 193.670 -30.250 194.080 -30.190 ;
        RECT 199.050 -29.890 199.460 -29.830 ;
        RECT 199.710 -29.890 200.860 -29.810 ;
        RECT 199.050 -30.190 200.860 -29.890 ;
        RECT 199.050 -30.250 199.460 -30.190 ;
        RECT 186.210 -30.370 186.660 -30.270 ;
        RECT 179.470 -31.520 179.910 -30.370 ;
        RECT 186.220 -31.520 186.660 -30.370 ;
        RECT 179.470 -32.170 180.620 -31.520 ;
        RECT 185.510 -32.170 186.660 -31.520 ;
        RECT 179.470 -33.320 179.910 -32.170 ;
        RECT 186.220 -33.320 186.660 -32.170 ;
        RECT 179.470 -33.420 179.920 -33.320 ;
        RECT 166.670 -33.500 167.080 -33.440 ;
        RECT 165.270 -33.800 167.080 -33.500 ;
        RECT 165.270 -33.880 166.420 -33.800 ;
        RECT 166.670 -33.860 167.080 -33.800 ;
        RECT 172.050 -33.500 172.460 -33.440 ;
        RECT 172.710 -33.500 173.860 -33.420 ;
        RECT 172.050 -33.800 173.860 -33.500 ;
        RECT 172.050 -33.860 172.460 -33.800 ;
        RECT 159.210 -33.980 159.660 -33.880 ;
        RECT 152.470 -35.130 152.910 -33.980 ;
        RECT 159.220 -35.130 159.660 -33.980 ;
        RECT 152.470 -35.780 153.620 -35.130 ;
        RECT 158.510 -35.780 159.660 -35.130 ;
        RECT 152.470 -36.930 152.910 -35.780 ;
        RECT 159.220 -36.930 159.660 -35.780 ;
        RECT 152.470 -37.030 152.920 -36.930 ;
        RECT 139.670 -37.110 140.080 -37.050 ;
        RECT 138.270 -37.410 140.080 -37.110 ;
        RECT 138.270 -37.490 139.420 -37.410 ;
        RECT 139.670 -37.470 140.080 -37.410 ;
        RECT 145.050 -37.110 145.460 -37.050 ;
        RECT 145.710 -37.110 146.860 -37.030 ;
        RECT 145.050 -37.410 146.860 -37.110 ;
        RECT 145.050 -37.470 145.460 -37.410 ;
        RECT 132.210 -37.590 132.660 -37.490 ;
        RECT 125.470 -38.740 125.910 -37.590 ;
        RECT 132.220 -38.740 132.660 -37.590 ;
        RECT 125.470 -39.390 126.620 -38.740 ;
        RECT 131.510 -39.390 132.660 -38.740 ;
        RECT 125.470 -40.540 125.910 -39.390 ;
        RECT 132.220 -40.540 132.660 -39.390 ;
        RECT 125.470 -40.640 125.920 -40.540 ;
        RECT 112.670 -40.720 113.080 -40.660 ;
        RECT 111.270 -40.940 113.080 -40.720 ;
        RECT 111.270 -41.090 111.720 -40.940 ;
        RECT 111.970 -40.980 113.080 -40.940 ;
        RECT 111.970 -41.090 112.420 -40.980 ;
        RECT 112.670 -41.080 113.080 -40.980 ;
        RECT 118.050 -40.720 118.460 -40.660 ;
        RECT 118.710 -40.720 119.860 -40.640 ;
        RECT 118.050 -40.940 119.860 -40.720 ;
        RECT 118.050 -40.980 119.160 -40.940 ;
        RECT 118.050 -41.080 118.460 -40.980 ;
        RECT 118.710 -41.090 119.160 -40.980 ;
        RECT 119.410 -41.090 119.860 -40.940 ;
        RECT 124.770 -40.720 125.920 -40.640 ;
        RECT 132.210 -40.640 132.660 -40.540 ;
        RECT 138.970 -37.590 139.420 -37.490 ;
        RECT 145.710 -37.490 146.860 -37.410 ;
        RECT 151.770 -37.110 152.920 -37.030 ;
        RECT 159.210 -37.030 159.660 -36.930 ;
        RECT 165.970 -33.980 166.420 -33.880 ;
        RECT 172.710 -33.880 173.860 -33.800 ;
        RECT 178.770 -33.500 179.920 -33.420 ;
        RECT 186.210 -33.420 186.660 -33.320 ;
        RECT 192.970 -30.370 193.420 -30.270 ;
        RECT 199.710 -30.270 200.860 -30.190 ;
        RECT 205.770 -29.890 206.920 -29.810 ;
        RECT 213.210 -29.810 213.660 -29.710 ;
        RECT 207.170 -29.890 207.580 -29.830 ;
        RECT 205.770 -30.190 207.580 -29.890 ;
        RECT 205.770 -30.270 206.920 -30.190 ;
        RECT 207.170 -30.250 207.580 -30.190 ;
        RECT 212.550 -29.890 212.960 -29.830 ;
        RECT 213.210 -29.890 214.360 -29.810 ;
        RECT 212.550 -30.190 214.360 -29.890 ;
        RECT 212.550 -30.250 212.960 -30.190 ;
        RECT 199.710 -30.370 200.160 -30.270 ;
        RECT 192.970 -31.520 193.410 -30.370 ;
        RECT 199.720 -31.520 200.160 -30.370 ;
        RECT 192.970 -32.170 194.120 -31.520 ;
        RECT 199.010 -32.170 200.160 -31.520 ;
        RECT 192.970 -33.320 193.410 -32.170 ;
        RECT 199.720 -33.320 200.160 -32.170 ;
        RECT 192.970 -33.420 193.420 -33.320 ;
        RECT 180.170 -33.500 180.580 -33.440 ;
        RECT 178.770 -33.800 180.580 -33.500 ;
        RECT 178.770 -33.880 179.920 -33.800 ;
        RECT 180.170 -33.860 180.580 -33.800 ;
        RECT 185.550 -33.500 185.960 -33.440 ;
        RECT 186.210 -33.500 187.360 -33.420 ;
        RECT 185.550 -33.800 187.360 -33.500 ;
        RECT 185.550 -33.860 185.960 -33.800 ;
        RECT 172.710 -33.980 173.160 -33.880 ;
        RECT 165.970 -35.130 166.410 -33.980 ;
        RECT 172.720 -35.130 173.160 -33.980 ;
        RECT 165.970 -35.780 167.120 -35.130 ;
        RECT 172.010 -35.780 173.160 -35.130 ;
        RECT 165.970 -36.930 166.410 -35.780 ;
        RECT 172.720 -36.930 173.160 -35.780 ;
        RECT 165.970 -37.030 166.420 -36.930 ;
        RECT 153.170 -37.110 153.580 -37.050 ;
        RECT 151.770 -37.410 153.580 -37.110 ;
        RECT 151.770 -37.490 152.920 -37.410 ;
        RECT 153.170 -37.470 153.580 -37.410 ;
        RECT 158.550 -37.110 158.960 -37.050 ;
        RECT 159.210 -37.110 160.360 -37.030 ;
        RECT 158.550 -37.410 160.360 -37.110 ;
        RECT 158.550 -37.470 158.960 -37.410 ;
        RECT 145.710 -37.590 146.160 -37.490 ;
        RECT 138.970 -38.740 139.410 -37.590 ;
        RECT 145.720 -38.740 146.160 -37.590 ;
        RECT 138.970 -39.390 140.120 -38.740 ;
        RECT 145.010 -39.390 146.160 -38.740 ;
        RECT 138.970 -40.540 139.410 -39.390 ;
        RECT 145.720 -40.540 146.160 -39.390 ;
        RECT 138.970 -40.640 139.420 -40.540 ;
        RECT 126.170 -40.720 126.580 -40.660 ;
        RECT 124.770 -40.940 126.580 -40.720 ;
        RECT 124.770 -41.090 125.220 -40.940 ;
        RECT 125.470 -40.980 126.580 -40.940 ;
        RECT 125.470 -41.090 125.920 -40.980 ;
        RECT 126.170 -41.080 126.580 -40.980 ;
        RECT 131.550 -40.720 131.960 -40.660 ;
        RECT 132.210 -40.720 133.360 -40.640 ;
        RECT 131.550 -40.940 133.360 -40.720 ;
        RECT 131.550 -40.980 132.660 -40.940 ;
        RECT 131.550 -41.080 131.960 -40.980 ;
        RECT 132.210 -41.090 132.660 -40.980 ;
        RECT 132.910 -41.090 133.360 -40.940 ;
        RECT 138.270 -40.720 139.420 -40.640 ;
        RECT 145.710 -40.640 146.160 -40.540 ;
        RECT 152.470 -37.590 152.920 -37.490 ;
        RECT 159.210 -37.490 160.360 -37.410 ;
        RECT 165.270 -37.110 166.420 -37.030 ;
        RECT 172.710 -37.030 173.160 -36.930 ;
        RECT 179.470 -33.980 179.920 -33.880 ;
        RECT 186.210 -33.880 187.360 -33.800 ;
        RECT 192.270 -33.500 193.420 -33.420 ;
        RECT 199.710 -33.420 200.160 -33.320 ;
        RECT 206.470 -30.370 206.920 -30.270 ;
        RECT 213.210 -30.270 214.360 -30.190 ;
        RECT 213.210 -30.370 213.660 -30.270 ;
        RECT 206.470 -31.520 206.910 -30.370 ;
        RECT 213.220 -31.520 213.660 -30.370 ;
        RECT 206.470 -32.170 207.620 -31.520 ;
        RECT 212.510 -32.170 213.660 -31.520 ;
        RECT 206.470 -33.320 206.910 -32.170 ;
        RECT 213.220 -33.320 213.660 -32.170 ;
        RECT 206.470 -33.420 206.920 -33.320 ;
        RECT 193.670 -33.500 194.080 -33.440 ;
        RECT 192.270 -33.800 194.080 -33.500 ;
        RECT 192.270 -33.880 193.420 -33.800 ;
        RECT 193.670 -33.860 194.080 -33.800 ;
        RECT 199.050 -33.500 199.460 -33.440 ;
        RECT 199.710 -33.500 200.860 -33.420 ;
        RECT 199.050 -33.800 200.860 -33.500 ;
        RECT 199.050 -33.860 199.460 -33.800 ;
        RECT 186.210 -33.980 186.660 -33.880 ;
        RECT 179.470 -35.130 179.910 -33.980 ;
        RECT 186.220 -35.130 186.660 -33.980 ;
        RECT 179.470 -35.780 180.620 -35.130 ;
        RECT 185.510 -35.780 186.660 -35.130 ;
        RECT 179.470 -36.930 179.910 -35.780 ;
        RECT 186.220 -36.930 186.660 -35.780 ;
        RECT 179.470 -37.030 179.920 -36.930 ;
        RECT 166.670 -37.110 167.080 -37.050 ;
        RECT 165.270 -37.410 167.080 -37.110 ;
        RECT 165.270 -37.490 166.420 -37.410 ;
        RECT 166.670 -37.470 167.080 -37.410 ;
        RECT 172.050 -37.110 172.460 -37.050 ;
        RECT 172.710 -37.110 173.860 -37.030 ;
        RECT 172.050 -37.410 173.860 -37.110 ;
        RECT 172.050 -37.470 172.460 -37.410 ;
        RECT 159.210 -37.590 159.660 -37.490 ;
        RECT 152.470 -38.740 152.910 -37.590 ;
        RECT 159.220 -38.740 159.660 -37.590 ;
        RECT 152.470 -39.390 153.620 -38.740 ;
        RECT 158.510 -39.390 159.660 -38.740 ;
        RECT 152.470 -40.540 152.910 -39.390 ;
        RECT 159.220 -40.540 159.660 -39.390 ;
        RECT 152.470 -40.640 152.920 -40.540 ;
        RECT 139.670 -40.720 140.080 -40.660 ;
        RECT 138.270 -40.940 140.080 -40.720 ;
        RECT 138.270 -41.090 138.720 -40.940 ;
        RECT 138.970 -40.980 140.080 -40.940 ;
        RECT 138.970 -41.090 139.420 -40.980 ;
        RECT 139.670 -41.080 140.080 -40.980 ;
        RECT 145.050 -40.720 145.460 -40.660 ;
        RECT 145.710 -40.720 146.860 -40.640 ;
        RECT 145.050 -40.940 146.860 -40.720 ;
        RECT 145.050 -40.980 146.160 -40.940 ;
        RECT 145.050 -41.080 145.460 -40.980 ;
        RECT 145.710 -41.090 146.160 -40.980 ;
        RECT 146.410 -41.090 146.860 -40.940 ;
        RECT 151.770 -40.720 152.920 -40.640 ;
        RECT 159.210 -40.640 159.660 -40.540 ;
        RECT 165.970 -37.590 166.420 -37.490 ;
        RECT 172.710 -37.490 173.860 -37.410 ;
        RECT 178.770 -37.110 179.920 -37.030 ;
        RECT 186.210 -37.030 186.660 -36.930 ;
        RECT 192.970 -33.980 193.420 -33.880 ;
        RECT 199.710 -33.880 200.860 -33.800 ;
        RECT 205.770 -33.500 206.920 -33.420 ;
        RECT 213.210 -33.420 213.660 -33.320 ;
        RECT 207.170 -33.500 207.580 -33.440 ;
        RECT 205.770 -33.800 207.580 -33.500 ;
        RECT 205.770 -33.880 206.920 -33.800 ;
        RECT 207.170 -33.860 207.580 -33.800 ;
        RECT 212.550 -33.500 212.960 -33.440 ;
        RECT 213.210 -33.500 214.360 -33.420 ;
        RECT 212.550 -33.800 214.360 -33.500 ;
        RECT 212.550 -33.860 212.960 -33.800 ;
        RECT 199.710 -33.980 200.160 -33.880 ;
        RECT 192.970 -35.130 193.410 -33.980 ;
        RECT 199.720 -35.130 200.160 -33.980 ;
        RECT 192.970 -35.780 194.120 -35.130 ;
        RECT 199.010 -35.780 200.160 -35.130 ;
        RECT 192.970 -36.930 193.410 -35.780 ;
        RECT 199.720 -36.930 200.160 -35.780 ;
        RECT 192.970 -37.030 193.420 -36.930 ;
        RECT 180.170 -37.110 180.580 -37.050 ;
        RECT 178.770 -37.410 180.580 -37.110 ;
        RECT 178.770 -37.490 179.920 -37.410 ;
        RECT 180.170 -37.470 180.580 -37.410 ;
        RECT 185.550 -37.110 185.960 -37.050 ;
        RECT 186.210 -37.110 187.360 -37.030 ;
        RECT 185.550 -37.410 187.360 -37.110 ;
        RECT 185.550 -37.470 185.960 -37.410 ;
        RECT 172.710 -37.590 173.160 -37.490 ;
        RECT 165.970 -38.740 166.410 -37.590 ;
        RECT 172.720 -38.740 173.160 -37.590 ;
        RECT 165.970 -39.390 167.120 -38.740 ;
        RECT 172.010 -39.390 173.160 -38.740 ;
        RECT 165.970 -40.540 166.410 -39.390 ;
        RECT 172.720 -40.540 173.160 -39.390 ;
        RECT 165.970 -40.640 166.420 -40.540 ;
        RECT 153.170 -40.720 153.580 -40.660 ;
        RECT 151.770 -40.940 153.580 -40.720 ;
        RECT 151.770 -41.090 152.220 -40.940 ;
        RECT 152.470 -40.980 153.580 -40.940 ;
        RECT 152.470 -41.090 152.920 -40.980 ;
        RECT 153.170 -41.080 153.580 -40.980 ;
        RECT 158.550 -40.720 158.960 -40.660 ;
        RECT 159.210 -40.720 160.360 -40.640 ;
        RECT 158.550 -40.940 160.360 -40.720 ;
        RECT 158.550 -40.980 159.660 -40.940 ;
        RECT 158.550 -41.080 158.960 -40.980 ;
        RECT 159.210 -41.090 159.660 -40.980 ;
        RECT 159.910 -41.090 160.360 -40.940 ;
        RECT 165.270 -40.720 166.420 -40.640 ;
        RECT 172.710 -40.640 173.160 -40.540 ;
        RECT 179.470 -37.590 179.920 -37.490 ;
        RECT 186.210 -37.490 187.360 -37.410 ;
        RECT 192.270 -37.110 193.420 -37.030 ;
        RECT 199.710 -37.030 200.160 -36.930 ;
        RECT 206.470 -33.980 206.920 -33.880 ;
        RECT 213.210 -33.880 214.360 -33.800 ;
        RECT 213.210 -33.980 213.660 -33.880 ;
        RECT 206.470 -35.130 206.910 -33.980 ;
        RECT 213.220 -35.130 213.660 -33.980 ;
        RECT 206.470 -35.780 207.620 -35.130 ;
        RECT 212.510 -35.780 213.660 -35.130 ;
        RECT 206.470 -36.930 206.910 -35.780 ;
        RECT 213.220 -36.930 213.660 -35.780 ;
        RECT 206.470 -37.030 206.920 -36.930 ;
        RECT 193.670 -37.110 194.080 -37.050 ;
        RECT 192.270 -37.410 194.080 -37.110 ;
        RECT 192.270 -37.490 193.420 -37.410 ;
        RECT 193.670 -37.470 194.080 -37.410 ;
        RECT 199.050 -37.110 199.460 -37.050 ;
        RECT 199.710 -37.110 200.860 -37.030 ;
        RECT 199.050 -37.410 200.860 -37.110 ;
        RECT 199.050 -37.470 199.460 -37.410 ;
        RECT 186.210 -37.590 186.660 -37.490 ;
        RECT 179.470 -38.740 179.910 -37.590 ;
        RECT 186.220 -38.740 186.660 -37.590 ;
        RECT 179.470 -39.390 180.620 -38.740 ;
        RECT 185.510 -39.390 186.660 -38.740 ;
        RECT 179.470 -40.540 179.910 -39.390 ;
        RECT 186.220 -40.540 186.660 -39.390 ;
        RECT 179.470 -40.640 179.920 -40.540 ;
        RECT 166.670 -40.720 167.080 -40.660 ;
        RECT 165.270 -40.940 167.080 -40.720 ;
        RECT 165.270 -41.090 165.720 -40.940 ;
        RECT 165.970 -40.980 167.080 -40.940 ;
        RECT 165.970 -41.090 166.420 -40.980 ;
        RECT 166.670 -41.080 167.080 -40.980 ;
        RECT 172.050 -40.720 172.460 -40.660 ;
        RECT 172.710 -40.720 173.860 -40.640 ;
        RECT 172.050 -40.940 173.860 -40.720 ;
        RECT 172.050 -40.980 173.160 -40.940 ;
        RECT 172.050 -41.080 172.460 -40.980 ;
        RECT 172.710 -41.090 173.160 -40.980 ;
        RECT 173.410 -41.090 173.860 -40.940 ;
        RECT 178.770 -40.720 179.920 -40.640 ;
        RECT 186.210 -40.640 186.660 -40.540 ;
        RECT 192.970 -37.590 193.420 -37.490 ;
        RECT 199.710 -37.490 200.860 -37.410 ;
        RECT 205.770 -37.110 206.920 -37.030 ;
        RECT 213.210 -37.030 213.660 -36.930 ;
        RECT 207.170 -37.110 207.580 -37.050 ;
        RECT 205.770 -37.410 207.580 -37.110 ;
        RECT 205.770 -37.490 206.920 -37.410 ;
        RECT 207.170 -37.470 207.580 -37.410 ;
        RECT 212.550 -37.110 212.960 -37.050 ;
        RECT 213.210 -37.110 214.360 -37.030 ;
        RECT 212.550 -37.410 214.360 -37.110 ;
        RECT 212.550 -37.470 212.960 -37.410 ;
        RECT 199.710 -37.590 200.160 -37.490 ;
        RECT 192.970 -38.740 193.410 -37.590 ;
        RECT 199.720 -38.740 200.160 -37.590 ;
        RECT 192.970 -39.390 194.120 -38.740 ;
        RECT 199.010 -39.390 200.160 -38.740 ;
        RECT 192.970 -40.540 193.410 -39.390 ;
        RECT 199.720 -40.540 200.160 -39.390 ;
        RECT 192.970 -40.640 193.420 -40.540 ;
        RECT 180.170 -40.720 180.580 -40.660 ;
        RECT 178.770 -40.940 180.580 -40.720 ;
        RECT 178.770 -41.090 179.220 -40.940 ;
        RECT 179.470 -40.980 180.580 -40.940 ;
        RECT 179.470 -41.090 179.920 -40.980 ;
        RECT 180.170 -41.080 180.580 -40.980 ;
        RECT 185.550 -40.720 185.960 -40.660 ;
        RECT 186.210 -40.720 187.360 -40.640 ;
        RECT 185.550 -40.940 187.360 -40.720 ;
        RECT 185.550 -40.980 186.660 -40.940 ;
        RECT 185.550 -41.080 185.960 -40.980 ;
        RECT 186.210 -41.090 186.660 -40.980 ;
        RECT 186.910 -41.090 187.360 -40.940 ;
        RECT 192.270 -40.720 193.420 -40.640 ;
        RECT 199.710 -40.640 200.160 -40.540 ;
        RECT 206.470 -37.590 206.920 -37.490 ;
        RECT 213.210 -37.490 214.360 -37.410 ;
        RECT 213.210 -37.590 213.660 -37.490 ;
        RECT 206.470 -38.740 206.910 -37.590 ;
        RECT 213.220 -38.740 213.660 -37.590 ;
        RECT 206.470 -39.390 207.620 -38.740 ;
        RECT 212.510 -39.390 213.660 -38.740 ;
        RECT 206.470 -40.540 206.910 -39.390 ;
        RECT 213.220 -40.540 213.660 -39.390 ;
        RECT 206.470 -40.640 206.920 -40.540 ;
        RECT 193.670 -40.720 194.080 -40.660 ;
        RECT 192.270 -40.940 194.080 -40.720 ;
        RECT 192.270 -41.090 192.720 -40.940 ;
        RECT 192.970 -40.980 194.080 -40.940 ;
        RECT 192.970 -41.090 193.420 -40.980 ;
        RECT 193.670 -41.080 194.080 -40.980 ;
        RECT 199.050 -40.720 199.460 -40.660 ;
        RECT 199.710 -40.720 200.860 -40.640 ;
        RECT 199.050 -40.940 200.860 -40.720 ;
        RECT 199.050 -40.980 200.160 -40.940 ;
        RECT 199.050 -41.080 199.460 -40.980 ;
        RECT 199.710 -41.090 200.160 -40.980 ;
        RECT 200.410 -41.090 200.860 -40.940 ;
        RECT 205.770 -40.720 206.920 -40.640 ;
        RECT 213.210 -40.640 213.660 -40.540 ;
        RECT 207.170 -40.720 207.580 -40.660 ;
        RECT 205.770 -40.940 207.580 -40.720 ;
        RECT 205.770 -41.090 206.220 -40.940 ;
        RECT 206.470 -40.980 207.580 -40.940 ;
        RECT 206.470 -41.090 206.920 -40.980 ;
        RECT 207.170 -41.080 207.580 -40.980 ;
        RECT 212.550 -40.720 212.960 -40.660 ;
        RECT 213.210 -40.720 214.360 -40.640 ;
        RECT 212.550 -40.940 214.360 -40.720 ;
        RECT 212.550 -40.980 213.660 -40.940 ;
        RECT 212.550 -41.080 212.960 -40.980 ;
        RECT 213.210 -41.090 213.660 -40.980 ;
        RECT 213.910 -41.090 214.360 -40.940 ;
      LAYER mcon ;
        RECT 4.050 16.760 4.310 17.020 ;
        RECT 10.820 16.760 11.080 17.020 ;
        RECT 17.550 16.760 17.810 17.020 ;
        RECT 24.320 16.760 24.580 17.020 ;
        RECT 4.060 14.950 4.310 15.220 ;
        RECT 10.820 14.950 11.070 15.220 ;
        RECT 31.050 16.760 31.310 17.020 ;
        RECT 37.820 16.760 38.080 17.020 ;
        RECT 17.560 14.950 17.810 15.220 ;
        RECT 24.320 14.950 24.570 15.220 ;
        RECT 4.050 13.150 4.310 13.410 ;
        RECT 10.820 13.150 11.080 13.410 ;
        RECT 44.550 16.760 44.810 17.020 ;
        RECT 51.320 16.760 51.580 17.020 ;
        RECT 31.060 14.950 31.310 15.220 ;
        RECT 37.820 14.950 38.070 15.220 ;
        RECT 17.550 13.150 17.810 13.410 ;
        RECT 24.320 13.150 24.580 13.410 ;
        RECT 4.060 11.340 4.310 11.610 ;
        RECT 10.820 11.340 11.070 11.610 ;
        RECT 58.050 16.760 58.310 17.020 ;
        RECT 64.820 16.760 65.080 17.020 ;
        RECT 44.560 14.950 44.810 15.220 ;
        RECT 51.320 14.950 51.570 15.220 ;
        RECT 31.050 13.150 31.310 13.410 ;
        RECT 37.820 13.150 38.080 13.410 ;
        RECT 17.560 11.340 17.810 11.610 ;
        RECT 24.320 11.340 24.570 11.610 ;
        RECT 4.050 9.540 4.310 9.800 ;
        RECT 10.820 9.540 11.080 9.800 ;
        RECT 71.550 16.760 71.810 17.020 ;
        RECT 78.320 16.760 78.580 17.020 ;
        RECT 58.060 14.950 58.310 15.220 ;
        RECT 64.820 14.950 65.070 15.220 ;
        RECT 44.550 13.150 44.810 13.410 ;
        RECT 51.320 13.150 51.580 13.410 ;
        RECT 31.060 11.340 31.310 11.610 ;
        RECT 37.820 11.340 38.070 11.610 ;
        RECT 17.550 9.540 17.810 9.800 ;
        RECT 24.320 9.540 24.580 9.800 ;
        RECT 4.060 7.730 4.310 8.000 ;
        RECT 10.820 7.730 11.070 8.000 ;
        RECT 85.050 16.760 85.310 17.020 ;
        RECT 91.820 16.760 92.080 17.020 ;
        RECT 71.560 14.950 71.810 15.220 ;
        RECT 78.320 14.950 78.570 15.220 ;
        RECT 58.050 13.150 58.310 13.410 ;
        RECT 64.820 13.150 65.080 13.410 ;
        RECT 44.560 11.340 44.810 11.610 ;
        RECT 51.320 11.340 51.570 11.610 ;
        RECT 31.050 9.540 31.310 9.800 ;
        RECT 37.820 9.540 38.080 9.800 ;
        RECT 17.560 7.730 17.810 8.000 ;
        RECT 24.320 7.730 24.570 8.000 ;
        RECT 4.050 5.930 4.310 6.190 ;
        RECT 10.820 5.930 11.080 6.190 ;
        RECT 98.550 16.760 98.810 17.020 ;
        RECT 105.320 16.760 105.580 17.020 ;
        RECT 85.060 14.950 85.310 15.220 ;
        RECT 91.820 14.950 92.070 15.220 ;
        RECT 71.550 13.150 71.810 13.410 ;
        RECT 78.320 13.150 78.580 13.410 ;
        RECT 58.060 11.340 58.310 11.610 ;
        RECT 64.820 11.340 65.070 11.610 ;
        RECT 44.550 9.540 44.810 9.800 ;
        RECT 51.320 9.540 51.580 9.800 ;
        RECT 31.060 7.730 31.310 8.000 ;
        RECT 37.820 7.730 38.070 8.000 ;
        RECT 17.550 5.930 17.810 6.190 ;
        RECT 24.320 5.930 24.580 6.190 ;
        RECT 4.060 4.120 4.310 4.390 ;
        RECT 10.820 4.120 11.070 4.390 ;
        RECT 112.050 16.760 112.310 17.020 ;
        RECT 118.820 16.760 119.080 17.020 ;
        RECT 98.560 14.950 98.810 15.220 ;
        RECT 105.320 14.950 105.570 15.220 ;
        RECT 85.050 13.150 85.310 13.410 ;
        RECT 91.820 13.150 92.080 13.410 ;
        RECT 71.560 11.340 71.810 11.610 ;
        RECT 78.320 11.340 78.570 11.610 ;
        RECT 58.050 9.540 58.310 9.800 ;
        RECT 64.820 9.540 65.080 9.800 ;
        RECT 44.560 7.730 44.810 8.000 ;
        RECT 51.320 7.730 51.570 8.000 ;
        RECT 31.050 5.930 31.310 6.190 ;
        RECT 37.820 5.930 38.080 6.190 ;
        RECT 17.560 4.120 17.810 4.390 ;
        RECT 24.320 4.120 24.570 4.390 ;
        RECT 4.050 2.320 4.310 2.580 ;
        RECT 10.820 2.320 11.080 2.580 ;
        RECT 125.550 16.760 125.810 17.020 ;
        RECT 132.320 16.760 132.580 17.020 ;
        RECT 112.060 14.950 112.310 15.220 ;
        RECT 118.820 14.950 119.070 15.220 ;
        RECT 98.550 13.150 98.810 13.410 ;
        RECT 105.320 13.150 105.580 13.410 ;
        RECT 85.060 11.340 85.310 11.610 ;
        RECT 91.820 11.340 92.070 11.610 ;
        RECT 71.550 9.540 71.810 9.800 ;
        RECT 78.320 9.540 78.580 9.800 ;
        RECT 58.060 7.730 58.310 8.000 ;
        RECT 64.820 7.730 65.070 8.000 ;
        RECT 44.550 5.930 44.810 6.190 ;
        RECT 51.320 5.930 51.580 6.190 ;
        RECT 31.060 4.120 31.310 4.390 ;
        RECT 37.820 4.120 38.070 4.390 ;
        RECT 17.550 2.320 17.810 2.580 ;
        RECT 24.320 2.320 24.580 2.580 ;
        RECT 4.060 0.510 4.310 0.780 ;
        RECT 10.820 0.510 11.070 0.780 ;
        RECT 139.050 16.760 139.310 17.020 ;
        RECT 145.820 16.760 146.080 17.020 ;
        RECT 125.560 14.950 125.810 15.220 ;
        RECT 132.320 14.950 132.570 15.220 ;
        RECT 112.050 13.150 112.310 13.410 ;
        RECT 118.820 13.150 119.080 13.410 ;
        RECT 98.560 11.340 98.810 11.610 ;
        RECT 105.320 11.340 105.570 11.610 ;
        RECT 85.050 9.540 85.310 9.800 ;
        RECT 91.820 9.540 92.080 9.800 ;
        RECT 71.560 7.730 71.810 8.000 ;
        RECT 78.320 7.730 78.570 8.000 ;
        RECT 58.050 5.930 58.310 6.190 ;
        RECT 64.820 5.930 65.080 6.190 ;
        RECT 44.560 4.120 44.810 4.390 ;
        RECT 51.320 4.120 51.570 4.390 ;
        RECT 31.050 2.320 31.310 2.580 ;
        RECT 37.820 2.320 38.080 2.580 ;
        RECT 17.560 0.510 17.810 0.780 ;
        RECT 24.320 0.510 24.570 0.780 ;
        RECT 4.050 -1.290 4.310 -1.030 ;
        RECT 10.820 -1.290 11.080 -1.030 ;
        RECT 152.550 16.760 152.810 17.020 ;
        RECT 159.320 16.760 159.580 17.020 ;
        RECT 139.060 14.950 139.310 15.220 ;
        RECT 145.820 14.950 146.070 15.220 ;
        RECT 125.550 13.150 125.810 13.410 ;
        RECT 132.320 13.150 132.580 13.410 ;
        RECT 112.060 11.340 112.310 11.610 ;
        RECT 118.820 11.340 119.070 11.610 ;
        RECT 98.550 9.540 98.810 9.800 ;
        RECT 105.320 9.540 105.580 9.800 ;
        RECT 85.060 7.730 85.310 8.000 ;
        RECT 91.820 7.730 92.070 8.000 ;
        RECT 71.550 5.930 71.810 6.190 ;
        RECT 78.320 5.930 78.580 6.190 ;
        RECT 58.060 4.120 58.310 4.390 ;
        RECT 64.820 4.120 65.070 4.390 ;
        RECT 44.550 2.320 44.810 2.580 ;
        RECT 51.320 2.320 51.580 2.580 ;
        RECT 31.060 0.510 31.310 0.780 ;
        RECT 37.820 0.510 38.070 0.780 ;
        RECT 17.550 -1.290 17.810 -1.030 ;
        RECT 24.320 -1.290 24.580 -1.030 ;
        RECT 4.060 -3.100 4.310 -2.830 ;
        RECT 10.820 -3.100 11.070 -2.830 ;
        RECT 166.050 16.760 166.310 17.020 ;
        RECT 172.820 16.760 173.080 17.020 ;
        RECT 152.560 14.950 152.810 15.220 ;
        RECT 159.320 14.950 159.570 15.220 ;
        RECT 139.050 13.150 139.310 13.410 ;
        RECT 145.820 13.150 146.080 13.410 ;
        RECT 125.560 11.340 125.810 11.610 ;
        RECT 132.320 11.340 132.570 11.610 ;
        RECT 112.050 9.540 112.310 9.800 ;
        RECT 118.820 9.540 119.080 9.800 ;
        RECT 98.560 7.730 98.810 8.000 ;
        RECT 105.320 7.730 105.570 8.000 ;
        RECT 85.050 5.930 85.310 6.190 ;
        RECT 91.820 5.930 92.080 6.190 ;
        RECT 71.560 4.120 71.810 4.390 ;
        RECT 78.320 4.120 78.570 4.390 ;
        RECT 58.050 2.320 58.310 2.580 ;
        RECT 64.820 2.320 65.080 2.580 ;
        RECT 44.560 0.510 44.810 0.780 ;
        RECT 51.320 0.510 51.570 0.780 ;
        RECT 31.050 -1.290 31.310 -1.030 ;
        RECT 37.820 -1.290 38.080 -1.030 ;
        RECT 17.560 -3.100 17.810 -2.830 ;
        RECT 24.320 -3.100 24.570 -2.830 ;
        RECT 4.050 -4.900 4.310 -4.640 ;
        RECT 10.820 -4.900 11.080 -4.640 ;
        RECT 179.550 16.760 179.810 17.020 ;
        RECT 186.320 16.760 186.580 17.020 ;
        RECT 166.060 14.950 166.310 15.220 ;
        RECT 172.820 14.950 173.070 15.220 ;
        RECT 152.550 13.150 152.810 13.410 ;
        RECT 159.320 13.150 159.580 13.410 ;
        RECT 139.060 11.340 139.310 11.610 ;
        RECT 145.820 11.340 146.070 11.610 ;
        RECT 125.550 9.540 125.810 9.800 ;
        RECT 132.320 9.540 132.580 9.800 ;
        RECT 112.060 7.730 112.310 8.000 ;
        RECT 118.820 7.730 119.070 8.000 ;
        RECT 98.550 5.930 98.810 6.190 ;
        RECT 105.320 5.930 105.580 6.190 ;
        RECT 85.060 4.120 85.310 4.390 ;
        RECT 91.820 4.120 92.070 4.390 ;
        RECT 71.550 2.320 71.810 2.580 ;
        RECT 78.320 2.320 78.580 2.580 ;
        RECT 58.060 0.510 58.310 0.780 ;
        RECT 64.820 0.510 65.070 0.780 ;
        RECT 44.550 -1.290 44.810 -1.030 ;
        RECT 51.320 -1.290 51.580 -1.030 ;
        RECT 31.060 -3.100 31.310 -2.830 ;
        RECT 37.820 -3.100 38.070 -2.830 ;
        RECT 17.550 -4.900 17.810 -4.640 ;
        RECT 24.320 -4.900 24.580 -4.640 ;
        RECT 4.060 -6.710 4.310 -6.440 ;
        RECT 10.820 -6.710 11.070 -6.440 ;
        RECT 193.050 16.760 193.310 17.020 ;
        RECT 199.820 16.760 200.080 17.020 ;
        RECT 179.560 14.950 179.810 15.220 ;
        RECT 186.320 14.950 186.570 15.220 ;
        RECT 166.050 13.150 166.310 13.410 ;
        RECT 172.820 13.150 173.080 13.410 ;
        RECT 152.560 11.340 152.810 11.610 ;
        RECT 159.320 11.340 159.570 11.610 ;
        RECT 139.050 9.540 139.310 9.800 ;
        RECT 145.820 9.540 146.080 9.800 ;
        RECT 125.560 7.730 125.810 8.000 ;
        RECT 132.320 7.730 132.570 8.000 ;
        RECT 112.050 5.930 112.310 6.190 ;
        RECT 118.820 5.930 119.080 6.190 ;
        RECT 98.560 4.120 98.810 4.390 ;
        RECT 105.320 4.120 105.570 4.390 ;
        RECT 85.050 2.320 85.310 2.580 ;
        RECT 91.820 2.320 92.080 2.580 ;
        RECT 71.560 0.510 71.810 0.780 ;
        RECT 78.320 0.510 78.570 0.780 ;
        RECT 58.050 -1.290 58.310 -1.030 ;
        RECT 64.820 -1.290 65.080 -1.030 ;
        RECT 44.560 -3.100 44.810 -2.830 ;
        RECT 51.320 -3.100 51.570 -2.830 ;
        RECT 31.050 -4.900 31.310 -4.640 ;
        RECT 37.820 -4.900 38.080 -4.640 ;
        RECT 17.560 -6.710 17.810 -6.440 ;
        RECT 24.320 -6.710 24.570 -6.440 ;
        RECT 4.050 -8.510 4.310 -8.250 ;
        RECT 10.820 -8.510 11.080 -8.250 ;
        RECT 206.550 16.760 206.810 17.020 ;
        RECT 213.320 16.760 213.580 17.020 ;
        RECT 193.060 14.950 193.310 15.220 ;
        RECT 199.820 14.950 200.070 15.220 ;
        RECT 179.550 13.150 179.810 13.410 ;
        RECT 186.320 13.150 186.580 13.410 ;
        RECT 166.060 11.340 166.310 11.610 ;
        RECT 172.820 11.340 173.070 11.610 ;
        RECT 152.550 9.540 152.810 9.800 ;
        RECT 159.320 9.540 159.580 9.800 ;
        RECT 139.060 7.730 139.310 8.000 ;
        RECT 145.820 7.730 146.070 8.000 ;
        RECT 125.550 5.930 125.810 6.190 ;
        RECT 132.320 5.930 132.580 6.190 ;
        RECT 112.060 4.120 112.310 4.390 ;
        RECT 118.820 4.120 119.070 4.390 ;
        RECT 98.550 2.320 98.810 2.580 ;
        RECT 105.320 2.320 105.580 2.580 ;
        RECT 85.060 0.510 85.310 0.780 ;
        RECT 91.820 0.510 92.070 0.780 ;
        RECT 71.550 -1.290 71.810 -1.030 ;
        RECT 78.320 -1.290 78.580 -1.030 ;
        RECT 58.060 -3.100 58.310 -2.830 ;
        RECT 64.820 -3.100 65.070 -2.830 ;
        RECT 44.550 -4.900 44.810 -4.640 ;
        RECT 51.320 -4.900 51.580 -4.640 ;
        RECT 31.060 -6.710 31.310 -6.440 ;
        RECT 37.820 -6.710 38.070 -6.440 ;
        RECT 17.550 -8.510 17.810 -8.250 ;
        RECT 24.320 -8.510 24.580 -8.250 ;
        RECT 4.060 -10.320 4.310 -10.050 ;
        RECT 10.820 -10.320 11.070 -10.050 ;
        RECT 206.560 14.950 206.810 15.220 ;
        RECT 213.320 14.950 213.570 15.220 ;
        RECT 193.050 13.150 193.310 13.410 ;
        RECT 199.820 13.150 200.080 13.410 ;
        RECT 179.560 11.340 179.810 11.610 ;
        RECT 186.320 11.340 186.570 11.610 ;
        RECT 166.050 9.540 166.310 9.800 ;
        RECT 172.820 9.540 173.080 9.800 ;
        RECT 152.560 7.730 152.810 8.000 ;
        RECT 159.320 7.730 159.570 8.000 ;
        RECT 139.050 5.930 139.310 6.190 ;
        RECT 145.820 5.930 146.080 6.190 ;
        RECT 125.560 4.120 125.810 4.390 ;
        RECT 132.320 4.120 132.570 4.390 ;
        RECT 112.050 2.320 112.310 2.580 ;
        RECT 118.820 2.320 119.080 2.580 ;
        RECT 98.560 0.510 98.810 0.780 ;
        RECT 105.320 0.510 105.570 0.780 ;
        RECT 85.050 -1.290 85.310 -1.030 ;
        RECT 91.820 -1.290 92.080 -1.030 ;
        RECT 71.560 -3.100 71.810 -2.830 ;
        RECT 78.320 -3.100 78.570 -2.830 ;
        RECT 58.050 -4.900 58.310 -4.640 ;
        RECT 64.820 -4.900 65.080 -4.640 ;
        RECT 44.560 -6.710 44.810 -6.440 ;
        RECT 51.320 -6.710 51.570 -6.440 ;
        RECT 31.050 -8.510 31.310 -8.250 ;
        RECT 37.820 -8.510 38.080 -8.250 ;
        RECT 17.560 -10.320 17.810 -10.050 ;
        RECT 24.320 -10.320 24.570 -10.050 ;
        RECT 4.050 -12.120 4.310 -11.860 ;
        RECT 10.820 -12.120 11.080 -11.860 ;
        RECT 206.550 13.150 206.810 13.410 ;
        RECT 213.320 13.150 213.580 13.410 ;
        RECT 193.060 11.340 193.310 11.610 ;
        RECT 199.820 11.340 200.070 11.610 ;
        RECT 179.550 9.540 179.810 9.800 ;
        RECT 186.320 9.540 186.580 9.800 ;
        RECT 166.060 7.730 166.310 8.000 ;
        RECT 172.820 7.730 173.070 8.000 ;
        RECT 152.550 5.930 152.810 6.190 ;
        RECT 159.320 5.930 159.580 6.190 ;
        RECT 139.060 4.120 139.310 4.390 ;
        RECT 145.820 4.120 146.070 4.390 ;
        RECT 125.550 2.320 125.810 2.580 ;
        RECT 132.320 2.320 132.580 2.580 ;
        RECT 112.060 0.510 112.310 0.780 ;
        RECT 118.820 0.510 119.070 0.780 ;
        RECT 98.550 -1.290 98.810 -1.030 ;
        RECT 105.320 -1.290 105.580 -1.030 ;
        RECT 85.060 -3.100 85.310 -2.830 ;
        RECT 91.820 -3.100 92.070 -2.830 ;
        RECT 71.550 -4.900 71.810 -4.640 ;
        RECT 78.320 -4.900 78.580 -4.640 ;
        RECT 58.060 -6.710 58.310 -6.440 ;
        RECT 64.820 -6.710 65.070 -6.440 ;
        RECT 44.550 -8.510 44.810 -8.250 ;
        RECT 51.320 -8.510 51.580 -8.250 ;
        RECT 31.060 -10.320 31.310 -10.050 ;
        RECT 37.820 -10.320 38.070 -10.050 ;
        RECT 17.550 -12.120 17.810 -11.860 ;
        RECT 24.320 -12.120 24.580 -11.860 ;
        RECT 4.060 -13.930 4.310 -13.660 ;
        RECT 10.820 -13.930 11.070 -13.660 ;
        RECT 206.560 11.340 206.810 11.610 ;
        RECT 213.320 11.340 213.570 11.610 ;
        RECT 193.050 9.540 193.310 9.800 ;
        RECT 199.820 9.540 200.080 9.800 ;
        RECT 179.560 7.730 179.810 8.000 ;
        RECT 186.320 7.730 186.570 8.000 ;
        RECT 166.050 5.930 166.310 6.190 ;
        RECT 172.820 5.930 173.080 6.190 ;
        RECT 152.560 4.120 152.810 4.390 ;
        RECT 159.320 4.120 159.570 4.390 ;
        RECT 139.050 2.320 139.310 2.580 ;
        RECT 145.820 2.320 146.080 2.580 ;
        RECT 125.560 0.510 125.810 0.780 ;
        RECT 132.320 0.510 132.570 0.780 ;
        RECT 112.050 -1.290 112.310 -1.030 ;
        RECT 118.820 -1.290 119.080 -1.030 ;
        RECT 98.560 -3.100 98.810 -2.830 ;
        RECT 105.320 -3.100 105.570 -2.830 ;
        RECT 85.050 -4.900 85.310 -4.640 ;
        RECT 91.820 -4.900 92.080 -4.640 ;
        RECT 71.560 -6.710 71.810 -6.440 ;
        RECT 78.320 -6.710 78.570 -6.440 ;
        RECT 58.050 -8.510 58.310 -8.250 ;
        RECT 64.820 -8.510 65.080 -8.250 ;
        RECT 44.560 -10.320 44.810 -10.050 ;
        RECT 51.320 -10.320 51.570 -10.050 ;
        RECT 31.050 -12.120 31.310 -11.860 ;
        RECT 37.820 -12.120 38.080 -11.860 ;
        RECT 17.560 -13.930 17.810 -13.660 ;
        RECT 24.320 -13.930 24.570 -13.660 ;
        RECT 4.050 -15.730 4.310 -15.470 ;
        RECT 10.820 -15.730 11.080 -15.470 ;
        RECT 206.550 9.540 206.810 9.800 ;
        RECT 213.320 9.540 213.580 9.800 ;
        RECT 193.060 7.730 193.310 8.000 ;
        RECT 199.820 7.730 200.070 8.000 ;
        RECT 179.550 5.930 179.810 6.190 ;
        RECT 186.320 5.930 186.580 6.190 ;
        RECT 166.060 4.120 166.310 4.390 ;
        RECT 172.820 4.120 173.070 4.390 ;
        RECT 152.550 2.320 152.810 2.580 ;
        RECT 159.320 2.320 159.580 2.580 ;
        RECT 139.060 0.510 139.310 0.780 ;
        RECT 145.820 0.510 146.070 0.780 ;
        RECT 125.550 -1.290 125.810 -1.030 ;
        RECT 132.320 -1.290 132.580 -1.030 ;
        RECT 112.060 -3.100 112.310 -2.830 ;
        RECT 118.820 -3.100 119.070 -2.830 ;
        RECT 98.550 -4.900 98.810 -4.640 ;
        RECT 105.320 -4.900 105.580 -4.640 ;
        RECT 85.060 -6.710 85.310 -6.440 ;
        RECT 91.820 -6.710 92.070 -6.440 ;
        RECT 71.550 -8.510 71.810 -8.250 ;
        RECT 78.320 -8.510 78.580 -8.250 ;
        RECT 58.060 -10.320 58.310 -10.050 ;
        RECT 64.820 -10.320 65.070 -10.050 ;
        RECT 44.550 -12.120 44.810 -11.860 ;
        RECT 51.320 -12.120 51.580 -11.860 ;
        RECT 31.060 -13.930 31.310 -13.660 ;
        RECT 37.820 -13.930 38.070 -13.660 ;
        RECT 17.550 -15.730 17.810 -15.470 ;
        RECT 24.320 -15.730 24.580 -15.470 ;
        RECT 4.060 -17.540 4.310 -17.270 ;
        RECT 10.820 -17.540 11.070 -17.270 ;
        RECT 206.560 7.730 206.810 8.000 ;
        RECT 213.320 7.730 213.570 8.000 ;
        RECT 193.050 5.930 193.310 6.190 ;
        RECT 199.820 5.930 200.080 6.190 ;
        RECT 179.560 4.120 179.810 4.390 ;
        RECT 186.320 4.120 186.570 4.390 ;
        RECT 166.050 2.320 166.310 2.580 ;
        RECT 172.820 2.320 173.080 2.580 ;
        RECT 152.560 0.510 152.810 0.780 ;
        RECT 159.320 0.510 159.570 0.780 ;
        RECT 139.050 -1.290 139.310 -1.030 ;
        RECT 145.820 -1.290 146.080 -1.030 ;
        RECT 125.560 -3.100 125.810 -2.830 ;
        RECT 132.320 -3.100 132.570 -2.830 ;
        RECT 112.050 -4.900 112.310 -4.640 ;
        RECT 118.820 -4.900 119.080 -4.640 ;
        RECT 98.560 -6.710 98.810 -6.440 ;
        RECT 105.320 -6.710 105.570 -6.440 ;
        RECT 85.050 -8.510 85.310 -8.250 ;
        RECT 91.820 -8.510 92.080 -8.250 ;
        RECT 71.560 -10.320 71.810 -10.050 ;
        RECT 78.320 -10.320 78.570 -10.050 ;
        RECT 58.050 -12.120 58.310 -11.860 ;
        RECT 64.820 -12.120 65.080 -11.860 ;
        RECT 44.560 -13.930 44.810 -13.660 ;
        RECT 51.320 -13.930 51.570 -13.660 ;
        RECT 31.050 -15.730 31.310 -15.470 ;
        RECT 37.820 -15.730 38.080 -15.470 ;
        RECT 17.560 -17.540 17.810 -17.270 ;
        RECT 24.320 -17.540 24.570 -17.270 ;
        RECT 4.050 -19.340 4.310 -19.080 ;
        RECT 10.820 -19.340 11.080 -19.080 ;
        RECT 206.550 5.930 206.810 6.190 ;
        RECT 213.320 5.930 213.580 6.190 ;
        RECT 193.060 4.120 193.310 4.390 ;
        RECT 199.820 4.120 200.070 4.390 ;
        RECT 179.550 2.320 179.810 2.580 ;
        RECT 186.320 2.320 186.580 2.580 ;
        RECT 166.060 0.510 166.310 0.780 ;
        RECT 172.820 0.510 173.070 0.780 ;
        RECT 152.550 -1.290 152.810 -1.030 ;
        RECT 159.320 -1.290 159.580 -1.030 ;
        RECT 139.060 -3.100 139.310 -2.830 ;
        RECT 145.820 -3.100 146.070 -2.830 ;
        RECT 125.550 -4.900 125.810 -4.640 ;
        RECT 132.320 -4.900 132.580 -4.640 ;
        RECT 112.060 -6.710 112.310 -6.440 ;
        RECT 118.820 -6.710 119.070 -6.440 ;
        RECT 98.550 -8.510 98.810 -8.250 ;
        RECT 105.320 -8.510 105.580 -8.250 ;
        RECT 85.060 -10.320 85.310 -10.050 ;
        RECT 91.820 -10.320 92.070 -10.050 ;
        RECT 71.550 -12.120 71.810 -11.860 ;
        RECT 78.320 -12.120 78.580 -11.860 ;
        RECT 58.060 -13.930 58.310 -13.660 ;
        RECT 64.820 -13.930 65.070 -13.660 ;
        RECT 44.550 -15.730 44.810 -15.470 ;
        RECT 51.320 -15.730 51.580 -15.470 ;
        RECT 31.060 -17.540 31.310 -17.270 ;
        RECT 37.820 -17.540 38.070 -17.270 ;
        RECT 17.550 -19.340 17.810 -19.080 ;
        RECT 24.320 -19.340 24.580 -19.080 ;
        RECT 4.060 -21.150 4.310 -20.880 ;
        RECT 10.820 -21.150 11.070 -20.880 ;
        RECT 206.560 4.120 206.810 4.390 ;
        RECT 213.320 4.120 213.570 4.390 ;
        RECT 193.050 2.320 193.310 2.580 ;
        RECT 199.820 2.320 200.080 2.580 ;
        RECT 179.560 0.510 179.810 0.780 ;
        RECT 186.320 0.510 186.570 0.780 ;
        RECT 166.050 -1.290 166.310 -1.030 ;
        RECT 172.820 -1.290 173.080 -1.030 ;
        RECT 152.560 -3.100 152.810 -2.830 ;
        RECT 159.320 -3.100 159.570 -2.830 ;
        RECT 139.050 -4.900 139.310 -4.640 ;
        RECT 145.820 -4.900 146.080 -4.640 ;
        RECT 125.560 -6.710 125.810 -6.440 ;
        RECT 132.320 -6.710 132.570 -6.440 ;
        RECT 112.050 -8.510 112.310 -8.250 ;
        RECT 118.820 -8.510 119.080 -8.250 ;
        RECT 98.560 -10.320 98.810 -10.050 ;
        RECT 105.320 -10.320 105.570 -10.050 ;
        RECT 85.050 -12.120 85.310 -11.860 ;
        RECT 91.820 -12.120 92.080 -11.860 ;
        RECT 71.560 -13.930 71.810 -13.660 ;
        RECT 78.320 -13.930 78.570 -13.660 ;
        RECT 58.050 -15.730 58.310 -15.470 ;
        RECT 64.820 -15.730 65.080 -15.470 ;
        RECT 44.560 -17.540 44.810 -17.270 ;
        RECT 51.320 -17.540 51.570 -17.270 ;
        RECT 31.050 -19.340 31.310 -19.080 ;
        RECT 37.820 -19.340 38.080 -19.080 ;
        RECT 17.560 -21.150 17.810 -20.880 ;
        RECT 24.320 -21.150 24.570 -20.880 ;
        RECT 4.050 -22.950 4.310 -22.690 ;
        RECT 10.820 -22.950 11.080 -22.690 ;
        RECT 206.550 2.320 206.810 2.580 ;
        RECT 213.320 2.320 213.580 2.580 ;
        RECT 193.060 0.510 193.310 0.780 ;
        RECT 199.820 0.510 200.070 0.780 ;
        RECT 179.550 -1.290 179.810 -1.030 ;
        RECT 186.320 -1.290 186.580 -1.030 ;
        RECT 166.060 -3.100 166.310 -2.830 ;
        RECT 172.820 -3.100 173.070 -2.830 ;
        RECT 152.550 -4.900 152.810 -4.640 ;
        RECT 159.320 -4.900 159.580 -4.640 ;
        RECT 139.060 -6.710 139.310 -6.440 ;
        RECT 145.820 -6.710 146.070 -6.440 ;
        RECT 125.550 -8.510 125.810 -8.250 ;
        RECT 132.320 -8.510 132.580 -8.250 ;
        RECT 112.060 -10.320 112.310 -10.050 ;
        RECT 118.820 -10.320 119.070 -10.050 ;
        RECT 98.550 -12.120 98.810 -11.860 ;
        RECT 105.320 -12.120 105.580 -11.860 ;
        RECT 85.060 -13.930 85.310 -13.660 ;
        RECT 91.820 -13.930 92.070 -13.660 ;
        RECT 71.550 -15.730 71.810 -15.470 ;
        RECT 78.320 -15.730 78.580 -15.470 ;
        RECT 58.060 -17.540 58.310 -17.270 ;
        RECT 64.820 -17.540 65.070 -17.270 ;
        RECT 44.550 -19.340 44.810 -19.080 ;
        RECT 51.320 -19.340 51.580 -19.080 ;
        RECT 31.060 -21.150 31.310 -20.880 ;
        RECT 37.820 -21.150 38.070 -20.880 ;
        RECT 17.550 -22.950 17.810 -22.690 ;
        RECT 24.320 -22.950 24.580 -22.690 ;
        RECT 4.060 -24.760 4.310 -24.490 ;
        RECT 10.820 -24.760 11.070 -24.490 ;
        RECT 206.560 0.510 206.810 0.780 ;
        RECT 213.320 0.510 213.570 0.780 ;
        RECT 193.050 -1.290 193.310 -1.030 ;
        RECT 199.820 -1.290 200.080 -1.030 ;
        RECT 179.560 -3.100 179.810 -2.830 ;
        RECT 186.320 -3.100 186.570 -2.830 ;
        RECT 166.050 -4.900 166.310 -4.640 ;
        RECT 172.820 -4.900 173.080 -4.640 ;
        RECT 152.560 -6.710 152.810 -6.440 ;
        RECT 159.320 -6.710 159.570 -6.440 ;
        RECT 139.050 -8.510 139.310 -8.250 ;
        RECT 145.820 -8.510 146.080 -8.250 ;
        RECT 125.560 -10.320 125.810 -10.050 ;
        RECT 132.320 -10.320 132.570 -10.050 ;
        RECT 112.050 -12.120 112.310 -11.860 ;
        RECT 118.820 -12.120 119.080 -11.860 ;
        RECT 98.560 -13.930 98.810 -13.660 ;
        RECT 105.320 -13.930 105.570 -13.660 ;
        RECT 85.050 -15.730 85.310 -15.470 ;
        RECT 91.820 -15.730 92.080 -15.470 ;
        RECT 71.560 -17.540 71.810 -17.270 ;
        RECT 78.320 -17.540 78.570 -17.270 ;
        RECT 58.050 -19.340 58.310 -19.080 ;
        RECT 64.820 -19.340 65.080 -19.080 ;
        RECT 44.560 -21.150 44.810 -20.880 ;
        RECT 51.320 -21.150 51.570 -20.880 ;
        RECT 31.050 -22.950 31.310 -22.690 ;
        RECT 37.820 -22.950 38.080 -22.690 ;
        RECT 17.560 -24.760 17.810 -24.490 ;
        RECT 24.320 -24.760 24.570 -24.490 ;
        RECT 4.050 -26.560 4.310 -26.300 ;
        RECT 10.820 -26.560 11.080 -26.300 ;
        RECT 206.550 -1.290 206.810 -1.030 ;
        RECT 213.320 -1.290 213.580 -1.030 ;
        RECT 193.060 -3.100 193.310 -2.830 ;
        RECT 199.820 -3.100 200.070 -2.830 ;
        RECT 179.550 -4.900 179.810 -4.640 ;
        RECT 186.320 -4.900 186.580 -4.640 ;
        RECT 166.060 -6.710 166.310 -6.440 ;
        RECT 172.820 -6.710 173.070 -6.440 ;
        RECT 152.550 -8.510 152.810 -8.250 ;
        RECT 159.320 -8.510 159.580 -8.250 ;
        RECT 139.060 -10.320 139.310 -10.050 ;
        RECT 145.820 -10.320 146.070 -10.050 ;
        RECT 125.550 -12.120 125.810 -11.860 ;
        RECT 132.320 -12.120 132.580 -11.860 ;
        RECT 112.060 -13.930 112.310 -13.660 ;
        RECT 118.820 -13.930 119.070 -13.660 ;
        RECT 98.550 -15.730 98.810 -15.470 ;
        RECT 105.320 -15.730 105.580 -15.470 ;
        RECT 85.060 -17.540 85.310 -17.270 ;
        RECT 91.820 -17.540 92.070 -17.270 ;
        RECT 71.550 -19.340 71.810 -19.080 ;
        RECT 78.320 -19.340 78.580 -19.080 ;
        RECT 58.060 -21.150 58.310 -20.880 ;
        RECT 64.820 -21.150 65.070 -20.880 ;
        RECT 44.550 -22.950 44.810 -22.690 ;
        RECT 51.320 -22.950 51.580 -22.690 ;
        RECT 31.060 -24.760 31.310 -24.490 ;
        RECT 37.820 -24.760 38.070 -24.490 ;
        RECT 17.550 -26.560 17.810 -26.300 ;
        RECT 24.320 -26.560 24.580 -26.300 ;
        RECT 4.060 -28.370 4.310 -28.100 ;
        RECT 10.820 -28.370 11.070 -28.100 ;
        RECT 206.560 -3.100 206.810 -2.830 ;
        RECT 213.320 -3.100 213.570 -2.830 ;
        RECT 193.050 -4.900 193.310 -4.640 ;
        RECT 199.820 -4.900 200.080 -4.640 ;
        RECT 179.560 -6.710 179.810 -6.440 ;
        RECT 186.320 -6.710 186.570 -6.440 ;
        RECT 166.050 -8.510 166.310 -8.250 ;
        RECT 172.820 -8.510 173.080 -8.250 ;
        RECT 152.560 -10.320 152.810 -10.050 ;
        RECT 159.320 -10.320 159.570 -10.050 ;
        RECT 139.050 -12.120 139.310 -11.860 ;
        RECT 145.820 -12.120 146.080 -11.860 ;
        RECT 125.560 -13.930 125.810 -13.660 ;
        RECT 132.320 -13.930 132.570 -13.660 ;
        RECT 112.050 -15.730 112.310 -15.470 ;
        RECT 118.820 -15.730 119.080 -15.470 ;
        RECT 98.560 -17.540 98.810 -17.270 ;
        RECT 105.320 -17.540 105.570 -17.270 ;
        RECT 85.050 -19.340 85.310 -19.080 ;
        RECT 91.820 -19.340 92.080 -19.080 ;
        RECT 71.560 -21.150 71.810 -20.880 ;
        RECT 78.320 -21.150 78.570 -20.880 ;
        RECT 58.050 -22.950 58.310 -22.690 ;
        RECT 64.820 -22.950 65.080 -22.690 ;
        RECT 44.560 -24.760 44.810 -24.490 ;
        RECT 51.320 -24.760 51.570 -24.490 ;
        RECT 31.050 -26.560 31.310 -26.300 ;
        RECT 37.820 -26.560 38.080 -26.300 ;
        RECT 17.560 -28.370 17.810 -28.100 ;
        RECT 24.320 -28.370 24.570 -28.100 ;
        RECT 4.050 -30.170 4.310 -29.910 ;
        RECT 10.820 -30.170 11.080 -29.910 ;
        RECT 206.550 -4.900 206.810 -4.640 ;
        RECT 213.320 -4.900 213.580 -4.640 ;
        RECT 193.060 -6.710 193.310 -6.440 ;
        RECT 199.820 -6.710 200.070 -6.440 ;
        RECT 179.550 -8.510 179.810 -8.250 ;
        RECT 186.320 -8.510 186.580 -8.250 ;
        RECT 166.060 -10.320 166.310 -10.050 ;
        RECT 172.820 -10.320 173.070 -10.050 ;
        RECT 152.550 -12.120 152.810 -11.860 ;
        RECT 159.320 -12.120 159.580 -11.860 ;
        RECT 139.060 -13.930 139.310 -13.660 ;
        RECT 145.820 -13.930 146.070 -13.660 ;
        RECT 125.550 -15.730 125.810 -15.470 ;
        RECT 132.320 -15.730 132.580 -15.470 ;
        RECT 112.060 -17.540 112.310 -17.270 ;
        RECT 118.820 -17.540 119.070 -17.270 ;
        RECT 98.550 -19.340 98.810 -19.080 ;
        RECT 105.320 -19.340 105.580 -19.080 ;
        RECT 85.060 -21.150 85.310 -20.880 ;
        RECT 91.820 -21.150 92.070 -20.880 ;
        RECT 71.550 -22.950 71.810 -22.690 ;
        RECT 78.320 -22.950 78.580 -22.690 ;
        RECT 58.060 -24.760 58.310 -24.490 ;
        RECT 64.820 -24.760 65.070 -24.490 ;
        RECT 44.550 -26.560 44.810 -26.300 ;
        RECT 51.320 -26.560 51.580 -26.300 ;
        RECT 31.060 -28.370 31.310 -28.100 ;
        RECT 37.820 -28.370 38.070 -28.100 ;
        RECT 17.550 -30.170 17.810 -29.910 ;
        RECT 24.320 -30.170 24.580 -29.910 ;
        RECT 4.060 -31.980 4.310 -31.710 ;
        RECT 10.820 -31.980 11.070 -31.710 ;
        RECT 206.560 -6.710 206.810 -6.440 ;
        RECT 213.320 -6.710 213.570 -6.440 ;
        RECT 193.050 -8.510 193.310 -8.250 ;
        RECT 199.820 -8.510 200.080 -8.250 ;
        RECT 179.560 -10.320 179.810 -10.050 ;
        RECT 186.320 -10.320 186.570 -10.050 ;
        RECT 166.050 -12.120 166.310 -11.860 ;
        RECT 172.820 -12.120 173.080 -11.860 ;
        RECT 152.560 -13.930 152.810 -13.660 ;
        RECT 159.320 -13.930 159.570 -13.660 ;
        RECT 139.050 -15.730 139.310 -15.470 ;
        RECT 145.820 -15.730 146.080 -15.470 ;
        RECT 125.560 -17.540 125.810 -17.270 ;
        RECT 132.320 -17.540 132.570 -17.270 ;
        RECT 112.050 -19.340 112.310 -19.080 ;
        RECT 118.820 -19.340 119.080 -19.080 ;
        RECT 98.560 -21.150 98.810 -20.880 ;
        RECT 105.320 -21.150 105.570 -20.880 ;
        RECT 85.050 -22.950 85.310 -22.690 ;
        RECT 91.820 -22.950 92.080 -22.690 ;
        RECT 71.560 -24.760 71.810 -24.490 ;
        RECT 78.320 -24.760 78.570 -24.490 ;
        RECT 58.050 -26.560 58.310 -26.300 ;
        RECT 64.820 -26.560 65.080 -26.300 ;
        RECT 44.560 -28.370 44.810 -28.100 ;
        RECT 51.320 -28.370 51.570 -28.100 ;
        RECT 31.050 -30.170 31.310 -29.910 ;
        RECT 37.820 -30.170 38.080 -29.910 ;
        RECT 17.560 -31.980 17.810 -31.710 ;
        RECT 24.320 -31.980 24.570 -31.710 ;
        RECT 4.050 -33.780 4.310 -33.520 ;
        RECT 10.820 -33.780 11.080 -33.520 ;
        RECT 206.550 -8.510 206.810 -8.250 ;
        RECT 213.320 -8.510 213.580 -8.250 ;
        RECT 193.060 -10.320 193.310 -10.050 ;
        RECT 199.820 -10.320 200.070 -10.050 ;
        RECT 179.550 -12.120 179.810 -11.860 ;
        RECT 186.320 -12.120 186.580 -11.860 ;
        RECT 166.060 -13.930 166.310 -13.660 ;
        RECT 172.820 -13.930 173.070 -13.660 ;
        RECT 152.550 -15.730 152.810 -15.470 ;
        RECT 159.320 -15.730 159.580 -15.470 ;
        RECT 139.060 -17.540 139.310 -17.270 ;
        RECT 145.820 -17.540 146.070 -17.270 ;
        RECT 125.550 -19.340 125.810 -19.080 ;
        RECT 132.320 -19.340 132.580 -19.080 ;
        RECT 112.060 -21.150 112.310 -20.880 ;
        RECT 118.820 -21.150 119.070 -20.880 ;
        RECT 98.550 -22.950 98.810 -22.690 ;
        RECT 105.320 -22.950 105.580 -22.690 ;
        RECT 85.060 -24.760 85.310 -24.490 ;
        RECT 91.820 -24.760 92.070 -24.490 ;
        RECT 71.550 -26.560 71.810 -26.300 ;
        RECT 78.320 -26.560 78.580 -26.300 ;
        RECT 58.060 -28.370 58.310 -28.100 ;
        RECT 64.820 -28.370 65.070 -28.100 ;
        RECT 44.550 -30.170 44.810 -29.910 ;
        RECT 51.320 -30.170 51.580 -29.910 ;
        RECT 31.060 -31.980 31.310 -31.710 ;
        RECT 37.820 -31.980 38.070 -31.710 ;
        RECT 17.550 -33.780 17.810 -33.520 ;
        RECT 24.320 -33.780 24.580 -33.520 ;
        RECT 4.060 -35.590 4.310 -35.320 ;
        RECT 10.820 -35.590 11.070 -35.320 ;
        RECT 206.560 -10.320 206.810 -10.050 ;
        RECT 213.320 -10.320 213.570 -10.050 ;
        RECT 193.050 -12.120 193.310 -11.860 ;
        RECT 199.820 -12.120 200.080 -11.860 ;
        RECT 179.560 -13.930 179.810 -13.660 ;
        RECT 186.320 -13.930 186.570 -13.660 ;
        RECT 166.050 -15.730 166.310 -15.470 ;
        RECT 172.820 -15.730 173.080 -15.470 ;
        RECT 152.560 -17.540 152.810 -17.270 ;
        RECT 159.320 -17.540 159.570 -17.270 ;
        RECT 139.050 -19.340 139.310 -19.080 ;
        RECT 145.820 -19.340 146.080 -19.080 ;
        RECT 125.560 -21.150 125.810 -20.880 ;
        RECT 132.320 -21.150 132.570 -20.880 ;
        RECT 112.050 -22.950 112.310 -22.690 ;
        RECT 118.820 -22.950 119.080 -22.690 ;
        RECT 98.560 -24.760 98.810 -24.490 ;
        RECT 105.320 -24.760 105.570 -24.490 ;
        RECT 85.050 -26.560 85.310 -26.300 ;
        RECT 91.820 -26.560 92.080 -26.300 ;
        RECT 71.560 -28.370 71.810 -28.100 ;
        RECT 78.320 -28.370 78.570 -28.100 ;
        RECT 58.050 -30.170 58.310 -29.910 ;
        RECT 64.820 -30.170 65.080 -29.910 ;
        RECT 44.560 -31.980 44.810 -31.710 ;
        RECT 51.320 -31.980 51.570 -31.710 ;
        RECT 31.050 -33.780 31.310 -33.520 ;
        RECT 37.820 -33.780 38.080 -33.520 ;
        RECT 17.560 -35.590 17.810 -35.320 ;
        RECT 24.320 -35.590 24.570 -35.320 ;
        RECT 4.050 -37.390 4.310 -37.130 ;
        RECT 10.820 -37.390 11.080 -37.130 ;
        RECT 206.550 -12.120 206.810 -11.860 ;
        RECT 213.320 -12.120 213.580 -11.860 ;
        RECT 193.060 -13.930 193.310 -13.660 ;
        RECT 199.820 -13.930 200.070 -13.660 ;
        RECT 179.550 -15.730 179.810 -15.470 ;
        RECT 186.320 -15.730 186.580 -15.470 ;
        RECT 166.060 -17.540 166.310 -17.270 ;
        RECT 172.820 -17.540 173.070 -17.270 ;
        RECT 152.550 -19.340 152.810 -19.080 ;
        RECT 159.320 -19.340 159.580 -19.080 ;
        RECT 139.060 -21.150 139.310 -20.880 ;
        RECT 145.820 -21.150 146.070 -20.880 ;
        RECT 125.550 -22.950 125.810 -22.690 ;
        RECT 132.320 -22.950 132.580 -22.690 ;
        RECT 112.060 -24.760 112.310 -24.490 ;
        RECT 118.820 -24.760 119.070 -24.490 ;
        RECT 98.550 -26.560 98.810 -26.300 ;
        RECT 105.320 -26.560 105.580 -26.300 ;
        RECT 85.060 -28.370 85.310 -28.100 ;
        RECT 91.820 -28.370 92.070 -28.100 ;
        RECT 71.550 -30.170 71.810 -29.910 ;
        RECT 78.320 -30.170 78.580 -29.910 ;
        RECT 58.060 -31.980 58.310 -31.710 ;
        RECT 64.820 -31.980 65.070 -31.710 ;
        RECT 44.550 -33.780 44.810 -33.520 ;
        RECT 51.320 -33.780 51.580 -33.520 ;
        RECT 31.060 -35.590 31.310 -35.320 ;
        RECT 37.820 -35.590 38.070 -35.320 ;
        RECT 17.550 -37.390 17.810 -37.130 ;
        RECT 24.320 -37.390 24.580 -37.130 ;
        RECT 4.060 -39.200 4.310 -38.930 ;
        RECT 10.820 -39.200 11.070 -38.930 ;
        RECT 206.560 -13.930 206.810 -13.660 ;
        RECT 213.320 -13.930 213.570 -13.660 ;
        RECT 193.050 -15.730 193.310 -15.470 ;
        RECT 199.820 -15.730 200.080 -15.470 ;
        RECT 179.560 -17.540 179.810 -17.270 ;
        RECT 186.320 -17.540 186.570 -17.270 ;
        RECT 166.050 -19.340 166.310 -19.080 ;
        RECT 172.820 -19.340 173.080 -19.080 ;
        RECT 152.560 -21.150 152.810 -20.880 ;
        RECT 159.320 -21.150 159.570 -20.880 ;
        RECT 139.050 -22.950 139.310 -22.690 ;
        RECT 145.820 -22.950 146.080 -22.690 ;
        RECT 125.560 -24.760 125.810 -24.490 ;
        RECT 132.320 -24.760 132.570 -24.490 ;
        RECT 112.050 -26.560 112.310 -26.300 ;
        RECT 118.820 -26.560 119.080 -26.300 ;
        RECT 98.560 -28.370 98.810 -28.100 ;
        RECT 105.320 -28.370 105.570 -28.100 ;
        RECT 85.050 -30.170 85.310 -29.910 ;
        RECT 91.820 -30.170 92.080 -29.910 ;
        RECT 71.560 -31.980 71.810 -31.710 ;
        RECT 78.320 -31.980 78.570 -31.710 ;
        RECT 58.050 -33.780 58.310 -33.520 ;
        RECT 64.820 -33.780 65.080 -33.520 ;
        RECT 44.560 -35.590 44.810 -35.320 ;
        RECT 51.320 -35.590 51.570 -35.320 ;
        RECT 31.050 -37.390 31.310 -37.130 ;
        RECT 37.820 -37.390 38.080 -37.130 ;
        RECT 17.560 -39.200 17.810 -38.930 ;
        RECT 24.320 -39.200 24.570 -38.930 ;
        RECT 4.050 -41.000 4.310 -40.740 ;
        RECT 10.820 -41.000 11.080 -40.740 ;
        RECT 206.550 -15.730 206.810 -15.470 ;
        RECT 213.320 -15.730 213.580 -15.470 ;
        RECT 193.060 -17.540 193.310 -17.270 ;
        RECT 199.820 -17.540 200.070 -17.270 ;
        RECT 179.550 -19.340 179.810 -19.080 ;
        RECT 186.320 -19.340 186.580 -19.080 ;
        RECT 166.060 -21.150 166.310 -20.880 ;
        RECT 172.820 -21.150 173.070 -20.880 ;
        RECT 152.550 -22.950 152.810 -22.690 ;
        RECT 159.320 -22.950 159.580 -22.690 ;
        RECT 139.060 -24.760 139.310 -24.490 ;
        RECT 145.820 -24.760 146.070 -24.490 ;
        RECT 125.550 -26.560 125.810 -26.300 ;
        RECT 132.320 -26.560 132.580 -26.300 ;
        RECT 112.060 -28.370 112.310 -28.100 ;
        RECT 118.820 -28.370 119.070 -28.100 ;
        RECT 98.550 -30.170 98.810 -29.910 ;
        RECT 105.320 -30.170 105.580 -29.910 ;
        RECT 85.060 -31.980 85.310 -31.710 ;
        RECT 91.820 -31.980 92.070 -31.710 ;
        RECT 71.550 -33.780 71.810 -33.520 ;
        RECT 78.320 -33.780 78.580 -33.520 ;
        RECT 58.060 -35.590 58.310 -35.320 ;
        RECT 64.820 -35.590 65.070 -35.320 ;
        RECT 44.550 -37.390 44.810 -37.130 ;
        RECT 51.320 -37.390 51.580 -37.130 ;
        RECT 31.060 -39.200 31.310 -38.930 ;
        RECT 37.820 -39.200 38.070 -38.930 ;
        RECT 17.550 -41.000 17.810 -40.740 ;
        RECT 24.320 -41.000 24.580 -40.740 ;
        RECT 206.560 -17.540 206.810 -17.270 ;
        RECT 213.320 -17.540 213.570 -17.270 ;
        RECT 193.050 -19.340 193.310 -19.080 ;
        RECT 199.820 -19.340 200.080 -19.080 ;
        RECT 179.560 -21.150 179.810 -20.880 ;
        RECT 186.320 -21.150 186.570 -20.880 ;
        RECT 166.050 -22.950 166.310 -22.690 ;
        RECT 172.820 -22.950 173.080 -22.690 ;
        RECT 152.560 -24.760 152.810 -24.490 ;
        RECT 159.320 -24.760 159.570 -24.490 ;
        RECT 139.050 -26.560 139.310 -26.300 ;
        RECT 145.820 -26.560 146.080 -26.300 ;
        RECT 125.560 -28.370 125.810 -28.100 ;
        RECT 132.320 -28.370 132.570 -28.100 ;
        RECT 112.050 -30.170 112.310 -29.910 ;
        RECT 118.820 -30.170 119.080 -29.910 ;
        RECT 98.560 -31.980 98.810 -31.710 ;
        RECT 105.320 -31.980 105.570 -31.710 ;
        RECT 85.050 -33.780 85.310 -33.520 ;
        RECT 91.820 -33.780 92.080 -33.520 ;
        RECT 71.560 -35.590 71.810 -35.320 ;
        RECT 78.320 -35.590 78.570 -35.320 ;
        RECT 58.050 -37.390 58.310 -37.130 ;
        RECT 64.820 -37.390 65.080 -37.130 ;
        RECT 44.560 -39.200 44.810 -38.930 ;
        RECT 51.320 -39.200 51.570 -38.930 ;
        RECT 31.050 -41.000 31.310 -40.740 ;
        RECT 37.820 -41.000 38.080 -40.740 ;
        RECT 206.550 -19.340 206.810 -19.080 ;
        RECT 213.320 -19.340 213.580 -19.080 ;
        RECT 193.060 -21.150 193.310 -20.880 ;
        RECT 199.820 -21.150 200.070 -20.880 ;
        RECT 179.550 -22.950 179.810 -22.690 ;
        RECT 186.320 -22.950 186.580 -22.690 ;
        RECT 166.060 -24.760 166.310 -24.490 ;
        RECT 172.820 -24.760 173.070 -24.490 ;
        RECT 152.550 -26.560 152.810 -26.300 ;
        RECT 159.320 -26.560 159.580 -26.300 ;
        RECT 139.060 -28.370 139.310 -28.100 ;
        RECT 145.820 -28.370 146.070 -28.100 ;
        RECT 125.550 -30.170 125.810 -29.910 ;
        RECT 132.320 -30.170 132.580 -29.910 ;
        RECT 112.060 -31.980 112.310 -31.710 ;
        RECT 118.820 -31.980 119.070 -31.710 ;
        RECT 98.550 -33.780 98.810 -33.520 ;
        RECT 105.320 -33.780 105.580 -33.520 ;
        RECT 85.060 -35.590 85.310 -35.320 ;
        RECT 91.820 -35.590 92.070 -35.320 ;
        RECT 71.550 -37.390 71.810 -37.130 ;
        RECT 78.320 -37.390 78.580 -37.130 ;
        RECT 58.060 -39.200 58.310 -38.930 ;
        RECT 64.820 -39.200 65.070 -38.930 ;
        RECT 44.550 -41.000 44.810 -40.740 ;
        RECT 51.320 -41.000 51.580 -40.740 ;
        RECT 206.560 -21.150 206.810 -20.880 ;
        RECT 213.320 -21.150 213.570 -20.880 ;
        RECT 193.050 -22.950 193.310 -22.690 ;
        RECT 199.820 -22.950 200.080 -22.690 ;
        RECT 179.560 -24.760 179.810 -24.490 ;
        RECT 186.320 -24.760 186.570 -24.490 ;
        RECT 166.050 -26.560 166.310 -26.300 ;
        RECT 172.820 -26.560 173.080 -26.300 ;
        RECT 152.560 -28.370 152.810 -28.100 ;
        RECT 159.320 -28.370 159.570 -28.100 ;
        RECT 139.050 -30.170 139.310 -29.910 ;
        RECT 145.820 -30.170 146.080 -29.910 ;
        RECT 125.560 -31.980 125.810 -31.710 ;
        RECT 132.320 -31.980 132.570 -31.710 ;
        RECT 112.050 -33.780 112.310 -33.520 ;
        RECT 118.820 -33.780 119.080 -33.520 ;
        RECT 98.560 -35.590 98.810 -35.320 ;
        RECT 105.320 -35.590 105.570 -35.320 ;
        RECT 85.050 -37.390 85.310 -37.130 ;
        RECT 91.820 -37.390 92.080 -37.130 ;
        RECT 71.560 -39.200 71.810 -38.930 ;
        RECT 78.320 -39.200 78.570 -38.930 ;
        RECT 58.050 -41.000 58.310 -40.740 ;
        RECT 64.820 -41.000 65.080 -40.740 ;
        RECT 206.550 -22.950 206.810 -22.690 ;
        RECT 213.320 -22.950 213.580 -22.690 ;
        RECT 193.060 -24.760 193.310 -24.490 ;
        RECT 199.820 -24.760 200.070 -24.490 ;
        RECT 179.550 -26.560 179.810 -26.300 ;
        RECT 186.320 -26.560 186.580 -26.300 ;
        RECT 166.060 -28.370 166.310 -28.100 ;
        RECT 172.820 -28.370 173.070 -28.100 ;
        RECT 152.550 -30.170 152.810 -29.910 ;
        RECT 159.320 -30.170 159.580 -29.910 ;
        RECT 139.060 -31.980 139.310 -31.710 ;
        RECT 145.820 -31.980 146.070 -31.710 ;
        RECT 125.550 -33.780 125.810 -33.520 ;
        RECT 132.320 -33.780 132.580 -33.520 ;
        RECT 112.060 -35.590 112.310 -35.320 ;
        RECT 118.820 -35.590 119.070 -35.320 ;
        RECT 98.550 -37.390 98.810 -37.130 ;
        RECT 105.320 -37.390 105.580 -37.130 ;
        RECT 85.060 -39.200 85.310 -38.930 ;
        RECT 91.820 -39.200 92.070 -38.930 ;
        RECT 71.550 -41.000 71.810 -40.740 ;
        RECT 78.320 -41.000 78.580 -40.740 ;
        RECT 206.560 -24.760 206.810 -24.490 ;
        RECT 213.320 -24.760 213.570 -24.490 ;
        RECT 193.050 -26.560 193.310 -26.300 ;
        RECT 199.820 -26.560 200.080 -26.300 ;
        RECT 179.560 -28.370 179.810 -28.100 ;
        RECT 186.320 -28.370 186.570 -28.100 ;
        RECT 166.050 -30.170 166.310 -29.910 ;
        RECT 172.820 -30.170 173.080 -29.910 ;
        RECT 152.560 -31.980 152.810 -31.710 ;
        RECT 159.320 -31.980 159.570 -31.710 ;
        RECT 139.050 -33.780 139.310 -33.520 ;
        RECT 145.820 -33.780 146.080 -33.520 ;
        RECT 125.560 -35.590 125.810 -35.320 ;
        RECT 132.320 -35.590 132.570 -35.320 ;
        RECT 112.050 -37.390 112.310 -37.130 ;
        RECT 118.820 -37.390 119.080 -37.130 ;
        RECT 98.560 -39.200 98.810 -38.930 ;
        RECT 105.320 -39.200 105.570 -38.930 ;
        RECT 85.050 -41.000 85.310 -40.740 ;
        RECT 91.820 -41.000 92.080 -40.740 ;
        RECT 206.550 -26.560 206.810 -26.300 ;
        RECT 213.320 -26.560 213.580 -26.300 ;
        RECT 193.060 -28.370 193.310 -28.100 ;
        RECT 199.820 -28.370 200.070 -28.100 ;
        RECT 179.550 -30.170 179.810 -29.910 ;
        RECT 186.320 -30.170 186.580 -29.910 ;
        RECT 166.060 -31.980 166.310 -31.710 ;
        RECT 172.820 -31.980 173.070 -31.710 ;
        RECT 152.550 -33.780 152.810 -33.520 ;
        RECT 159.320 -33.780 159.580 -33.520 ;
        RECT 139.060 -35.590 139.310 -35.320 ;
        RECT 145.820 -35.590 146.070 -35.320 ;
        RECT 125.550 -37.390 125.810 -37.130 ;
        RECT 132.320 -37.390 132.580 -37.130 ;
        RECT 112.060 -39.200 112.310 -38.930 ;
        RECT 118.820 -39.200 119.070 -38.930 ;
        RECT 98.550 -41.000 98.810 -40.740 ;
        RECT 105.320 -41.000 105.580 -40.740 ;
        RECT 206.560 -28.370 206.810 -28.100 ;
        RECT 213.320 -28.370 213.570 -28.100 ;
        RECT 193.050 -30.170 193.310 -29.910 ;
        RECT 199.820 -30.170 200.080 -29.910 ;
        RECT 179.560 -31.980 179.810 -31.710 ;
        RECT 186.320 -31.980 186.570 -31.710 ;
        RECT 166.050 -33.780 166.310 -33.520 ;
        RECT 172.820 -33.780 173.080 -33.520 ;
        RECT 152.560 -35.590 152.810 -35.320 ;
        RECT 159.320 -35.590 159.570 -35.320 ;
        RECT 139.050 -37.390 139.310 -37.130 ;
        RECT 145.820 -37.390 146.080 -37.130 ;
        RECT 125.560 -39.200 125.810 -38.930 ;
        RECT 132.320 -39.200 132.570 -38.930 ;
        RECT 112.050 -41.000 112.310 -40.740 ;
        RECT 118.820 -41.000 119.080 -40.740 ;
        RECT 206.550 -30.170 206.810 -29.910 ;
        RECT 213.320 -30.170 213.580 -29.910 ;
        RECT 193.060 -31.980 193.310 -31.710 ;
        RECT 199.820 -31.980 200.070 -31.710 ;
        RECT 179.550 -33.780 179.810 -33.520 ;
        RECT 186.320 -33.780 186.580 -33.520 ;
        RECT 166.060 -35.590 166.310 -35.320 ;
        RECT 172.820 -35.590 173.070 -35.320 ;
        RECT 152.550 -37.390 152.810 -37.130 ;
        RECT 159.320 -37.390 159.580 -37.130 ;
        RECT 139.060 -39.200 139.310 -38.930 ;
        RECT 145.820 -39.200 146.070 -38.930 ;
        RECT 125.550 -41.000 125.810 -40.740 ;
        RECT 132.320 -41.000 132.580 -40.740 ;
        RECT 206.560 -31.980 206.810 -31.710 ;
        RECT 213.320 -31.980 213.570 -31.710 ;
        RECT 193.050 -33.780 193.310 -33.520 ;
        RECT 199.820 -33.780 200.080 -33.520 ;
        RECT 179.560 -35.590 179.810 -35.320 ;
        RECT 186.320 -35.590 186.570 -35.320 ;
        RECT 166.050 -37.390 166.310 -37.130 ;
        RECT 172.820 -37.390 173.080 -37.130 ;
        RECT 152.560 -39.200 152.810 -38.930 ;
        RECT 159.320 -39.200 159.570 -38.930 ;
        RECT 139.050 -41.000 139.310 -40.740 ;
        RECT 145.820 -41.000 146.080 -40.740 ;
        RECT 206.550 -33.780 206.810 -33.520 ;
        RECT 213.320 -33.780 213.580 -33.520 ;
        RECT 193.060 -35.590 193.310 -35.320 ;
        RECT 199.820 -35.590 200.070 -35.320 ;
        RECT 179.550 -37.390 179.810 -37.130 ;
        RECT 186.320 -37.390 186.580 -37.130 ;
        RECT 166.060 -39.200 166.310 -38.930 ;
        RECT 172.820 -39.200 173.070 -38.930 ;
        RECT 152.550 -41.000 152.810 -40.740 ;
        RECT 159.320 -41.000 159.580 -40.740 ;
        RECT 206.560 -35.590 206.810 -35.320 ;
        RECT 213.320 -35.590 213.570 -35.320 ;
        RECT 193.050 -37.390 193.310 -37.130 ;
        RECT 199.820 -37.390 200.080 -37.130 ;
        RECT 179.560 -39.200 179.810 -38.930 ;
        RECT 186.320 -39.200 186.570 -38.930 ;
        RECT 166.050 -41.000 166.310 -40.740 ;
        RECT 172.820 -41.000 173.080 -40.740 ;
        RECT 206.550 -37.390 206.810 -37.130 ;
        RECT 213.320 -37.390 213.580 -37.130 ;
        RECT 193.060 -39.200 193.310 -38.930 ;
        RECT 199.820 -39.200 200.070 -38.930 ;
        RECT 179.550 -41.000 179.810 -40.740 ;
        RECT 186.320 -41.000 186.580 -40.740 ;
        RECT 206.560 -39.200 206.810 -38.930 ;
        RECT 213.320 -39.200 213.570 -38.930 ;
        RECT 193.050 -41.000 193.310 -40.740 ;
        RECT 199.820 -41.000 200.080 -40.740 ;
        RECT 206.550 -41.000 206.810 -40.740 ;
        RECT 213.320 -41.000 213.580 -40.740 ;
      LAYER met1 ;
        RECT 3.920 -43.310 4.470 19.330 ;
        RECT 10.660 -43.350 11.210 19.370 ;
        RECT 17.420 -43.350 17.970 19.370 ;
        RECT 24.160 -43.350 24.710 19.370 ;
        RECT 30.920 -43.350 31.470 19.370 ;
        RECT 37.660 -43.350 38.210 19.370 ;
        RECT 44.420 -43.350 44.970 19.370 ;
        RECT 51.160 -43.310 51.710 19.330 ;
        RECT 57.920 -43.310 58.470 19.330 ;
        RECT 64.660 -43.350 65.210 19.370 ;
        RECT 71.420 -43.350 71.970 19.370 ;
        RECT 78.160 -43.350 78.710 19.370 ;
        RECT 84.920 -43.350 85.470 19.370 ;
        RECT 91.660 -43.350 92.210 19.370 ;
        RECT 98.420 -43.350 98.970 19.370 ;
        RECT 105.160 -43.310 105.710 19.330 ;
        RECT 111.920 -43.310 112.470 19.330 ;
        RECT 118.660 -43.350 119.210 19.370 ;
        RECT 125.420 -43.350 125.970 19.370 ;
        RECT 132.160 -43.350 132.710 19.370 ;
        RECT 138.920 -43.350 139.470 19.370 ;
        RECT 145.660 -43.350 146.210 19.370 ;
        RECT 152.420 -43.350 152.970 19.370 ;
        RECT 159.160 -43.310 159.710 19.330 ;
        RECT 165.920 -43.310 166.470 19.330 ;
        RECT 172.660 -43.350 173.210 19.370 ;
        RECT 179.420 -43.350 179.970 19.370 ;
        RECT 186.160 -43.350 186.710 19.370 ;
        RECT 192.920 -43.350 193.470 19.370 ;
        RECT 199.660 -43.350 200.210 19.370 ;
        RECT 206.420 -43.350 206.970 19.370 ;
        RECT 213.160 -43.310 213.710 19.330 ;
      LAYER via ;
        RECT 4.020 18.270 4.380 18.610 ;
        RECT 10.760 18.250 11.120 18.590 ;
        RECT 17.490 18.350 17.850 18.690 ;
        RECT 24.280 18.350 24.640 18.690 ;
        RECT 31.040 18.310 31.400 18.650 ;
        RECT 37.800 18.280 38.160 18.620 ;
        RECT 44.530 18.220 44.890 18.560 ;
        RECT 51.230 18.220 51.590 18.560 ;
        RECT 58.010 18.240 58.370 18.580 ;
        RECT 64.760 18.270 65.120 18.610 ;
        RECT 71.560 18.250 71.920 18.590 ;
        RECT 78.270 18.240 78.630 18.580 ;
        RECT 85.010 18.260 85.370 18.600 ;
        RECT 91.730 18.210 92.090 18.550 ;
        RECT 98.520 18.210 98.880 18.550 ;
        RECT 105.280 18.240 105.640 18.580 ;
        RECT 112.000 18.180 112.360 18.520 ;
        RECT 118.790 18.170 119.150 18.510 ;
        RECT 125.490 18.230 125.850 18.570 ;
        RECT 132.280 18.310 132.640 18.650 ;
        RECT 139.040 18.350 139.400 18.690 ;
        RECT 145.790 18.320 146.150 18.660 ;
        RECT 152.520 18.290 152.880 18.630 ;
        RECT 159.240 18.280 159.600 18.620 ;
        RECT 166.030 18.380 166.390 18.720 ;
        RECT 172.740 18.380 173.100 18.720 ;
        RECT 179.500 18.380 179.860 18.720 ;
        RECT 186.280 18.370 186.640 18.710 ;
        RECT 193.020 18.360 193.380 18.700 ;
        RECT 199.780 18.290 200.140 18.630 ;
        RECT 206.530 18.290 206.890 18.630 ;
        RECT 213.240 18.280 213.600 18.620 ;
      LAYER met2 ;
        RECT -0.790 17.920 221.150 18.980 ;
    END
  END vccd1
  PIN vssd1
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.600 17.070 1.040 17.110 ;
        RECT -0.060 17.020 1.040 17.070 ;
        RECT 1.420 17.020 1.870 17.120 ;
        RECT -0.060 16.770 1.870 17.020 ;
        RECT -0.060 16.750 1.040 16.770 ;
        RECT 0.600 16.680 1.040 16.750 ;
        RECT 1.420 16.760 1.870 16.770 ;
        RECT 1.420 16.550 2.950 16.760 ;
        RECT 2.500 16.270 2.950 16.550 ;
        RECT 2.500 13.620 2.950 13.900 ;
        RECT 0.600 13.410 1.040 13.500 ;
        RECT 1.420 13.410 2.950 13.620 ;
        RECT 0.600 13.400 1.870 13.410 ;
        RECT 0.390 13.210 1.870 13.400 ;
        RECT 0.600 13.150 1.870 13.210 ;
        RECT 0.600 13.060 1.040 13.150 ;
        RECT 1.420 12.940 2.950 13.150 ;
        RECT 2.500 12.660 2.950 12.940 ;
        RECT 2.500 10.010 2.950 10.290 ;
        RECT 0.600 9.800 1.040 9.890 ;
        RECT 1.420 9.800 2.950 10.010 ;
        RECT 0.600 9.540 1.870 9.800 ;
        RECT 0.600 9.450 1.040 9.540 ;
        RECT 1.420 9.330 2.950 9.540 ;
        RECT 2.500 9.050 2.950 9.330 ;
        RECT 2.500 6.400 2.950 6.680 ;
        RECT 0.600 6.190 1.040 6.280 ;
        RECT 1.420 6.190 2.950 6.400 ;
        RECT 0.600 6.130 1.870 6.190 ;
        RECT 0.390 5.940 1.870 6.130 ;
        RECT 0.600 5.930 1.870 5.940 ;
        RECT 0.600 5.840 1.040 5.930 ;
        RECT 1.420 5.720 2.950 5.930 ;
        RECT 2.500 5.440 2.950 5.720 ;
        RECT 2.500 2.790 2.950 3.070 ;
        RECT 0.600 2.630 1.040 2.670 ;
        RECT -0.060 2.580 1.040 2.630 ;
        RECT 1.420 2.580 2.950 2.790 ;
        RECT -0.060 2.320 1.870 2.580 ;
        RECT -0.060 2.270 1.040 2.320 ;
        RECT 0.600 2.230 1.040 2.270 ;
        RECT 1.420 2.110 2.950 2.320 ;
        RECT 2.500 1.830 2.950 2.110 ;
        RECT 2.500 -0.820 2.950 -0.540 ;
        RECT 0.600 -1.030 1.040 -0.940 ;
        RECT 1.420 -1.030 2.950 -0.820 ;
        RECT 0.600 -1.040 1.870 -1.030 ;
        RECT 0.390 -1.230 1.870 -1.040 ;
        RECT 0.600 -1.290 1.870 -1.230 ;
        RECT 0.600 -1.380 1.040 -1.290 ;
        RECT 1.420 -1.500 2.950 -1.290 ;
        RECT 2.500 -1.780 2.950 -1.500 ;
        RECT 2.500 -4.430 2.950 -4.150 ;
        RECT 0.600 -4.640 1.040 -4.550 ;
        RECT 1.420 -4.640 2.950 -4.430 ;
        RECT 0.600 -4.900 1.870 -4.640 ;
        RECT 0.600 -4.990 1.040 -4.900 ;
        RECT 1.420 -5.110 2.950 -4.900 ;
        RECT 2.500 -5.390 2.950 -5.110 ;
        RECT 2.500 -8.040 2.950 -7.760 ;
        RECT 0.600 -8.250 1.040 -8.160 ;
        RECT 1.420 -8.250 2.950 -8.040 ;
        RECT 0.600 -8.310 1.870 -8.250 ;
        RECT 0.390 -8.500 1.870 -8.310 ;
        RECT 0.600 -8.510 1.870 -8.500 ;
        RECT 0.600 -8.600 1.040 -8.510 ;
        RECT 1.420 -8.720 2.950 -8.510 ;
        RECT 2.500 -9.000 2.950 -8.720 ;
        RECT 2.500 -11.650 2.950 -11.370 ;
        RECT 0.600 -11.810 1.040 -11.770 ;
        RECT -0.060 -11.860 1.040 -11.810 ;
        RECT 1.420 -11.860 2.950 -11.650 ;
        RECT -0.060 -12.120 1.870 -11.860 ;
        RECT -0.060 -12.170 1.040 -12.120 ;
        RECT 0.600 -12.210 1.040 -12.170 ;
        RECT 1.420 -12.330 2.950 -12.120 ;
        RECT 2.500 -12.610 2.950 -12.330 ;
        RECT 2.500 -15.260 2.950 -14.980 ;
        RECT 0.600 -15.470 1.040 -15.380 ;
        RECT 1.420 -15.470 2.950 -15.260 ;
        RECT 0.600 -15.480 1.870 -15.470 ;
        RECT 0.390 -15.670 1.870 -15.480 ;
        RECT 0.600 -15.730 1.870 -15.670 ;
        RECT 0.600 -15.820 1.040 -15.730 ;
        RECT 1.420 -15.940 2.950 -15.730 ;
        RECT 2.500 -16.220 2.950 -15.940 ;
        RECT 2.500 -18.870 2.950 -18.590 ;
        RECT 0.600 -19.080 1.040 -18.990 ;
        RECT 1.420 -19.080 2.950 -18.870 ;
        RECT 0.600 -19.340 1.870 -19.080 ;
        RECT 0.600 -19.430 1.040 -19.340 ;
        RECT 1.420 -19.550 2.950 -19.340 ;
        RECT 2.500 -19.830 2.950 -19.550 ;
        RECT 2.500 -22.480 2.950 -22.200 ;
        RECT 0.600 -22.690 1.040 -22.600 ;
        RECT 1.420 -22.690 2.950 -22.480 ;
        RECT 0.600 -22.750 1.870 -22.690 ;
        RECT 0.390 -22.940 1.870 -22.750 ;
        RECT 0.600 -22.950 1.870 -22.940 ;
        RECT 0.600 -23.040 1.040 -22.950 ;
        RECT 1.420 -23.160 2.950 -22.950 ;
        RECT 2.500 -23.440 2.950 -23.160 ;
        RECT 2.500 -26.090 2.950 -25.810 ;
        RECT 0.600 -26.250 1.040 -26.210 ;
        RECT -0.060 -26.300 1.040 -26.250 ;
        RECT 1.420 -26.300 2.950 -26.090 ;
        RECT -0.060 -26.560 1.870 -26.300 ;
        RECT -0.060 -26.610 1.040 -26.560 ;
        RECT 0.600 -26.650 1.040 -26.610 ;
        RECT 1.420 -26.770 2.950 -26.560 ;
        RECT 2.500 -27.050 2.950 -26.770 ;
        RECT 2.500 -29.700 2.950 -29.420 ;
        RECT 0.600 -29.910 1.040 -29.820 ;
        RECT 1.420 -29.910 2.950 -29.700 ;
        RECT 0.600 -29.920 1.870 -29.910 ;
        RECT 0.390 -30.110 1.870 -29.920 ;
        RECT 0.600 -30.170 1.870 -30.110 ;
        RECT 0.600 -30.260 1.040 -30.170 ;
        RECT 1.420 -30.380 2.950 -30.170 ;
        RECT 2.500 -30.660 2.950 -30.380 ;
        RECT 2.500 -33.310 2.950 -33.030 ;
        RECT 0.600 -33.520 1.040 -33.430 ;
        RECT 1.420 -33.520 2.950 -33.310 ;
        RECT 0.600 -33.780 1.870 -33.520 ;
        RECT 0.600 -33.870 1.040 -33.780 ;
        RECT 1.420 -33.990 2.950 -33.780 ;
        RECT 2.500 -34.270 2.950 -33.990 ;
        RECT 2.500 -36.920 2.950 -36.640 ;
        RECT 0.600 -37.130 1.040 -37.040 ;
        RECT 1.420 -37.130 2.950 -36.920 ;
        RECT 0.600 -37.190 1.870 -37.130 ;
        RECT 0.390 -37.380 1.870 -37.190 ;
        RECT 0.600 -37.390 1.870 -37.380 ;
        RECT 0.600 -37.480 1.040 -37.390 ;
        RECT 1.420 -37.600 2.950 -37.390 ;
        RECT 2.500 -37.880 2.950 -37.600 ;
        RECT 2.500 -40.530 2.950 -40.250 ;
        RECT 0.600 -40.730 1.040 -40.660 ;
        RECT -0.060 -40.750 1.040 -40.730 ;
        RECT 1.420 -40.740 2.950 -40.530 ;
        RECT 1.420 -40.750 1.870 -40.740 ;
        RECT -0.060 -41.000 1.870 -40.750 ;
        RECT -0.060 -41.050 1.040 -41.000 ;
        RECT 0.600 -41.090 1.040 -41.050 ;
        RECT 1.420 -41.100 1.870 -41.000 ;
      LAYER mcon ;
        RECT 2.600 16.370 2.860 16.630 ;
        RECT 2.600 13.540 2.860 13.800 ;
        RECT 2.600 12.760 2.860 13.020 ;
        RECT 2.600 9.930 2.860 10.190 ;
        RECT 2.600 9.150 2.860 9.410 ;
        RECT 2.600 6.320 2.860 6.580 ;
        RECT 2.600 5.540 2.860 5.800 ;
        RECT 2.600 2.710 2.860 2.970 ;
        RECT 2.600 1.930 2.860 2.190 ;
        RECT 2.600 -0.900 2.860 -0.640 ;
        RECT 2.600 -1.680 2.860 -1.420 ;
        RECT 2.600 -4.510 2.860 -4.250 ;
        RECT 2.600 -5.290 2.860 -5.030 ;
        RECT 2.600 -8.120 2.860 -7.860 ;
        RECT 2.600 -8.900 2.860 -8.640 ;
        RECT 2.600 -11.730 2.860 -11.470 ;
        RECT 2.600 -12.510 2.860 -12.250 ;
        RECT 2.600 -15.340 2.860 -15.080 ;
        RECT 2.600 -16.120 2.860 -15.860 ;
        RECT 2.600 -18.950 2.860 -18.690 ;
        RECT 2.600 -19.730 2.860 -19.470 ;
        RECT 2.600 -22.560 2.860 -22.300 ;
        RECT 2.600 -23.340 2.860 -23.080 ;
        RECT 2.600 -26.170 2.860 -25.910 ;
        RECT 2.600 -26.950 2.860 -26.690 ;
        RECT 2.600 -29.780 2.860 -29.520 ;
        RECT 2.600 -30.560 2.860 -30.300 ;
        RECT 2.600 -33.390 2.860 -33.130 ;
        RECT 2.600 -34.170 2.860 -33.910 ;
        RECT 2.600 -37.000 2.860 -36.740 ;
        RECT 2.600 -37.780 2.860 -37.520 ;
        RECT 2.600 -40.610 2.860 -40.350 ;
      LAYER met1 ;
        RECT 2.500 -41.200 3.070 17.220 ;
        RECT 5.360 -41.220 5.950 17.240 ;
      LAYER via ;
        RECT 2.650 15.130 2.910 15.390 ;
        RECT 2.650 14.780 2.910 15.040 ;
        RECT 2.650 11.520 2.910 11.780 ;
        RECT 2.650 11.170 2.910 11.430 ;
        RECT 2.650 7.910 2.910 8.170 ;
        RECT 2.650 7.560 2.910 7.820 ;
        RECT 2.650 4.300 2.910 4.560 ;
        RECT 2.650 3.950 2.910 4.210 ;
        RECT 2.650 0.690 2.910 0.950 ;
        RECT 2.650 0.340 2.910 0.600 ;
        RECT 2.650 -2.920 2.910 -2.660 ;
        RECT 2.650 -3.270 2.910 -3.010 ;
        RECT 2.650 -6.530 2.910 -6.270 ;
        RECT 2.650 -6.880 2.910 -6.620 ;
        RECT 2.650 -10.140 2.910 -9.880 ;
        RECT 2.650 -10.490 2.910 -10.230 ;
        RECT 2.650 -13.750 2.910 -13.490 ;
        RECT 2.650 -14.100 2.910 -13.840 ;
        RECT 2.650 -17.360 2.910 -17.100 ;
        RECT 2.650 -17.710 2.910 -17.450 ;
        RECT 2.650 -20.970 2.910 -20.710 ;
        RECT 2.650 -21.320 2.910 -21.060 ;
        RECT 2.650 -24.580 2.910 -24.320 ;
        RECT 2.650 -24.930 2.910 -24.670 ;
        RECT 2.650 -28.190 2.910 -27.930 ;
        RECT 2.650 -28.540 2.910 -28.280 ;
        RECT 2.650 -31.800 2.910 -31.540 ;
        RECT 2.650 -32.150 2.910 -31.890 ;
        RECT 2.650 -35.410 2.910 -35.150 ;
        RECT 2.650 -35.760 2.910 -35.500 ;
        RECT 2.650 -39.020 2.910 -38.760 ;
        RECT 2.650 -39.370 2.910 -39.110 ;
        RECT 5.510 15.140 5.770 15.400 ;
        RECT 5.510 14.770 5.770 15.030 ;
        RECT 5.510 11.530 5.770 11.790 ;
        RECT 5.510 11.160 5.770 11.420 ;
        RECT 5.510 7.920 5.770 8.180 ;
        RECT 5.510 7.550 5.770 7.810 ;
        RECT 5.510 4.310 5.770 4.570 ;
        RECT 5.510 3.940 5.770 4.200 ;
        RECT 5.510 0.700 5.770 0.960 ;
        RECT 5.510 0.330 5.770 0.590 ;
        RECT 5.510 -2.910 5.770 -2.650 ;
        RECT 5.510 -3.280 5.770 -3.020 ;
        RECT 5.510 -6.520 5.770 -6.260 ;
        RECT 5.510 -6.890 5.770 -6.630 ;
        RECT 5.510 -10.130 5.770 -9.870 ;
        RECT 5.510 -10.500 5.770 -10.240 ;
        RECT 5.510 -13.740 5.770 -13.480 ;
        RECT 5.510 -14.110 5.770 -13.850 ;
        RECT 5.510 -17.350 5.770 -17.090 ;
        RECT 5.510 -17.720 5.770 -17.460 ;
        RECT 5.510 -20.960 5.770 -20.700 ;
        RECT 5.510 -21.330 5.770 -21.070 ;
        RECT 5.510 -24.570 5.770 -24.310 ;
        RECT 5.510 -24.940 5.770 -24.680 ;
        RECT 5.510 -28.180 5.770 -27.920 ;
        RECT 5.510 -28.550 5.770 -28.290 ;
        RECT 5.510 -31.790 5.770 -31.530 ;
        RECT 5.510 -32.160 5.770 -31.900 ;
        RECT 5.510 -35.400 5.770 -35.140 ;
        RECT 5.510 -35.770 5.770 -35.510 ;
        RECT 5.510 -39.010 5.770 -38.750 ;
        RECT 5.510 -39.380 5.770 -39.120 ;
      LAYER met2 ;
        RECT 2.560 15.410 3.020 15.490 ;
        RECT 5.420 15.410 5.870 15.500 ;
        RECT 2.560 15.180 5.870 15.410 ;
        RECT 2.560 14.990 3.020 15.180 ;
        RECT 5.420 14.990 5.870 15.180 ;
        RECT 2.560 14.760 5.870 14.990 ;
        RECT 2.560 14.680 3.020 14.760 ;
        RECT 5.420 14.670 5.870 14.760 ;
        RECT 2.560 11.800 3.020 11.880 ;
        RECT 5.420 11.800 5.870 11.890 ;
        RECT 2.560 11.570 5.870 11.800 ;
        RECT 2.560 11.380 3.020 11.570 ;
        RECT 5.420 11.380 5.870 11.570 ;
        RECT 2.560 11.150 5.870 11.380 ;
        RECT 2.560 11.070 3.020 11.150 ;
        RECT 5.420 11.060 5.870 11.150 ;
        RECT 2.560 8.190 3.020 8.270 ;
        RECT 5.420 8.190 5.870 8.280 ;
        RECT 2.560 7.960 5.870 8.190 ;
        RECT 2.560 7.770 3.020 7.960 ;
        RECT 5.420 7.770 5.870 7.960 ;
        RECT 2.560 7.540 5.870 7.770 ;
        RECT 2.560 7.460 3.020 7.540 ;
        RECT 5.420 7.450 5.870 7.540 ;
        RECT 2.560 4.580 3.020 4.660 ;
        RECT 5.420 4.580 5.870 4.670 ;
        RECT 2.560 4.350 5.870 4.580 ;
        RECT 2.560 4.160 3.020 4.350 ;
        RECT 5.420 4.160 5.870 4.350 ;
        RECT 2.560 3.930 5.870 4.160 ;
        RECT 2.560 3.850 3.020 3.930 ;
        RECT 5.420 3.840 5.870 3.930 ;
        RECT 2.560 0.970 3.020 1.050 ;
        RECT 5.420 0.970 5.870 1.060 ;
        RECT 2.560 0.740 5.870 0.970 ;
        RECT 2.560 0.550 3.020 0.740 ;
        RECT 5.420 0.550 5.870 0.740 ;
        RECT 2.560 0.320 5.870 0.550 ;
        RECT 2.560 0.240 3.020 0.320 ;
        RECT 5.420 0.230 5.870 0.320 ;
        RECT 2.560 -2.640 3.020 -2.560 ;
        RECT 5.420 -2.640 5.870 -2.550 ;
        RECT 2.560 -2.870 5.870 -2.640 ;
        RECT 2.560 -3.060 3.020 -2.870 ;
        RECT 5.420 -3.060 5.870 -2.870 ;
        RECT 2.560 -3.290 5.870 -3.060 ;
        RECT 2.560 -3.370 3.020 -3.290 ;
        RECT 5.420 -3.380 5.870 -3.290 ;
        RECT 2.560 -6.250 3.020 -6.170 ;
        RECT 5.420 -6.250 5.870 -6.160 ;
        RECT 2.560 -6.480 5.870 -6.250 ;
        RECT 2.560 -6.670 3.020 -6.480 ;
        RECT 5.420 -6.670 5.870 -6.480 ;
        RECT 2.560 -6.900 5.870 -6.670 ;
        RECT 2.560 -6.980 3.020 -6.900 ;
        RECT 5.420 -6.990 5.870 -6.900 ;
        RECT 2.560 -9.860 3.020 -9.780 ;
        RECT 5.420 -9.860 5.870 -9.770 ;
        RECT 2.560 -10.090 5.870 -9.860 ;
        RECT 2.560 -10.280 3.020 -10.090 ;
        RECT 5.420 -10.280 5.870 -10.090 ;
        RECT 2.560 -10.510 5.870 -10.280 ;
        RECT 2.560 -10.590 3.020 -10.510 ;
        RECT 5.420 -10.600 5.870 -10.510 ;
        RECT 2.560 -13.470 3.020 -13.390 ;
        RECT 5.420 -13.470 5.870 -13.380 ;
        RECT 2.560 -13.700 5.870 -13.470 ;
        RECT 2.560 -13.890 3.020 -13.700 ;
        RECT 5.420 -13.890 5.870 -13.700 ;
        RECT 2.560 -14.120 5.870 -13.890 ;
        RECT 2.560 -14.200 3.020 -14.120 ;
        RECT 5.420 -14.210 5.870 -14.120 ;
        RECT 2.560 -17.080 3.020 -17.000 ;
        RECT 5.420 -17.080 5.870 -16.990 ;
        RECT 2.560 -17.310 5.870 -17.080 ;
        RECT 2.560 -17.500 3.020 -17.310 ;
        RECT 5.420 -17.500 5.870 -17.310 ;
        RECT 2.560 -17.730 5.870 -17.500 ;
        RECT 2.560 -17.810 3.020 -17.730 ;
        RECT 5.420 -17.820 5.870 -17.730 ;
        RECT 2.560 -20.690 3.020 -20.610 ;
        RECT 5.420 -20.690 5.870 -20.600 ;
        RECT 2.560 -20.920 5.870 -20.690 ;
        RECT 2.560 -21.110 3.020 -20.920 ;
        RECT 5.420 -21.110 5.870 -20.920 ;
        RECT 2.560 -21.340 5.870 -21.110 ;
        RECT 2.560 -21.420 3.020 -21.340 ;
        RECT 5.420 -21.430 5.870 -21.340 ;
        RECT 2.560 -24.300 3.020 -24.220 ;
        RECT 5.420 -24.300 5.870 -24.210 ;
        RECT 2.560 -24.530 5.870 -24.300 ;
        RECT 2.560 -24.720 3.020 -24.530 ;
        RECT 5.420 -24.720 5.870 -24.530 ;
        RECT 2.560 -24.950 5.870 -24.720 ;
        RECT 2.560 -25.030 3.020 -24.950 ;
        RECT 5.420 -25.040 5.870 -24.950 ;
        RECT 2.560 -27.910 3.020 -27.830 ;
        RECT 5.420 -27.910 5.870 -27.820 ;
        RECT 2.560 -28.140 5.870 -27.910 ;
        RECT 2.560 -28.330 3.020 -28.140 ;
        RECT 5.420 -28.330 5.870 -28.140 ;
        RECT 2.560 -28.560 5.870 -28.330 ;
        RECT 2.560 -28.640 3.020 -28.560 ;
        RECT 5.420 -28.650 5.870 -28.560 ;
        RECT 2.560 -31.520 3.020 -31.440 ;
        RECT 5.420 -31.520 5.870 -31.430 ;
        RECT 2.560 -31.750 5.870 -31.520 ;
        RECT 2.560 -31.940 3.020 -31.750 ;
        RECT 5.420 -31.940 5.870 -31.750 ;
        RECT 2.560 -32.170 5.870 -31.940 ;
        RECT 2.560 -32.250 3.020 -32.170 ;
        RECT 5.420 -32.260 5.870 -32.170 ;
        RECT 2.560 -35.130 3.020 -35.050 ;
        RECT 5.420 -35.130 5.870 -35.040 ;
        RECT 2.560 -35.360 5.870 -35.130 ;
        RECT 2.560 -35.550 3.020 -35.360 ;
        RECT 5.420 -35.550 5.870 -35.360 ;
        RECT 2.560 -35.780 5.870 -35.550 ;
        RECT 2.560 -35.860 3.020 -35.780 ;
        RECT 5.420 -35.870 5.870 -35.780 ;
        RECT 2.560 -38.740 3.020 -38.660 ;
        RECT 5.420 -38.740 5.870 -38.650 ;
        RECT 2.560 -38.970 5.870 -38.740 ;
        RECT 2.560 -39.160 3.020 -38.970 ;
        RECT 5.420 -39.160 5.870 -38.970 ;
        RECT 2.560 -39.390 5.870 -39.160 ;
        RECT 2.560 -39.470 3.020 -39.390 ;
        RECT 5.420 -39.480 5.870 -39.390 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 13.260 17.020 13.710 17.120 ;
        RECT 14.090 17.020 14.540 17.110 ;
        RECT 14.920 17.020 15.370 17.120 ;
        RECT 13.260 16.770 15.370 17.020 ;
        RECT 13.260 16.760 13.710 16.770 ;
        RECT 12.180 16.550 13.710 16.760 ;
        RECT 14.090 16.680 14.540 16.770 ;
        RECT 14.920 16.760 15.370 16.770 ;
        RECT 26.760 17.020 27.210 17.120 ;
        RECT 27.590 17.020 28.040 17.110 ;
        RECT 28.420 17.020 28.870 17.120 ;
        RECT 26.760 16.770 28.870 17.020 ;
        RECT 26.760 16.760 27.210 16.770 ;
        RECT 14.920 16.550 16.450 16.760 ;
        RECT 1.420 16.100 1.870 16.210 ;
        RECT 3.270 16.100 3.720 16.210 ;
        RECT 1.420 15.860 3.720 16.100 ;
        RECT 1.420 15.760 1.870 15.860 ;
        RECT 2.260 15.430 2.670 15.860 ;
        RECT 3.270 15.790 3.720 15.860 ;
        RECT 4.670 16.100 5.120 16.180 ;
        RECT 5.720 16.100 6.130 16.540 ;
        RECT 6.520 16.100 6.970 16.210 ;
        RECT 4.670 15.860 6.970 16.100 ;
        RECT 4.670 15.760 5.120 15.860 ;
        RECT 6.520 15.760 6.970 15.860 ;
        RECT 8.160 16.100 8.610 16.210 ;
        RECT 9.000 16.100 9.410 16.540 ;
        RECT 12.180 16.270 12.630 16.550 ;
        RECT 16.000 16.270 16.450 16.550 ;
        RECT 25.680 16.550 27.210 16.760 ;
        RECT 27.590 16.680 28.040 16.770 ;
        RECT 28.420 16.760 28.870 16.770 ;
        RECT 40.260 17.020 40.710 17.120 ;
        RECT 41.090 17.020 41.540 17.110 ;
        RECT 41.920 17.020 42.370 17.120 ;
        RECT 40.260 16.770 42.370 17.020 ;
        RECT 40.260 16.760 40.710 16.770 ;
        RECT 28.420 16.550 29.950 16.760 ;
        RECT 10.010 16.100 10.460 16.180 ;
        RECT 8.160 15.860 10.460 16.100 ;
        RECT 8.160 15.760 8.610 15.860 ;
        RECT 10.010 15.760 10.460 15.860 ;
        RECT 11.410 16.100 11.860 16.210 ;
        RECT 13.260 16.100 13.710 16.210 ;
        RECT 11.410 15.860 13.710 16.100 ;
        RECT 11.410 15.790 11.860 15.860 ;
        RECT 5.420 15.280 6.970 15.500 ;
        RECT 5.420 14.890 5.920 15.280 ;
        RECT 6.520 15.230 6.970 15.280 ;
        RECT 7.350 15.230 7.780 15.290 ;
        RECT 8.160 15.280 9.710 15.500 ;
        RECT 12.460 15.430 12.870 15.860 ;
        RECT 13.260 15.760 13.710 15.860 ;
        RECT 14.920 16.100 15.370 16.210 ;
        RECT 16.770 16.100 17.220 16.210 ;
        RECT 14.920 15.860 17.220 16.100 ;
        RECT 14.920 15.760 15.370 15.860 ;
        RECT 15.760 15.430 16.170 15.860 ;
        RECT 16.770 15.790 17.220 15.860 ;
        RECT 18.170 16.100 18.620 16.180 ;
        RECT 19.220 16.100 19.630 16.540 ;
        RECT 20.020 16.100 20.470 16.210 ;
        RECT 18.170 15.860 20.470 16.100 ;
        RECT 18.170 15.760 18.620 15.860 ;
        RECT 20.020 15.760 20.470 15.860 ;
        RECT 21.660 16.100 22.110 16.210 ;
        RECT 22.500 16.100 22.910 16.540 ;
        RECT 25.680 16.270 26.130 16.550 ;
        RECT 29.500 16.270 29.950 16.550 ;
        RECT 39.180 16.550 40.710 16.760 ;
        RECT 41.090 16.680 41.540 16.770 ;
        RECT 41.920 16.760 42.370 16.770 ;
        RECT 53.760 17.070 54.210 17.120 ;
        RECT 54.590 17.070 55.040 17.110 ;
        RECT 55.420 17.070 55.870 17.120 ;
        RECT 53.760 16.760 55.870 17.070 ;
        RECT 67.260 17.020 67.710 17.120 ;
        RECT 68.090 17.020 68.540 17.110 ;
        RECT 68.920 17.020 69.370 17.120 ;
        RECT 67.260 16.770 69.370 17.020 ;
        RECT 67.260 16.760 67.710 16.770 ;
        RECT 41.920 16.550 43.450 16.760 ;
        RECT 23.510 16.100 23.960 16.180 ;
        RECT 21.660 15.860 23.960 16.100 ;
        RECT 21.660 15.760 22.110 15.860 ;
        RECT 23.510 15.760 23.960 15.860 ;
        RECT 24.910 16.100 25.360 16.210 ;
        RECT 26.760 16.100 27.210 16.210 ;
        RECT 24.910 15.860 27.210 16.100 ;
        RECT 24.910 15.790 25.360 15.860 ;
        RECT 8.160 15.230 8.610 15.280 ;
        RECT 6.520 14.940 8.610 15.230 ;
        RECT 6.520 14.890 6.970 14.940 ;
        RECT 1.420 14.310 1.870 14.410 ;
        RECT 2.260 14.310 2.670 14.740 ;
        RECT 5.420 14.670 6.970 14.890 ;
        RECT 7.350 14.880 7.780 14.940 ;
        RECT 8.160 14.890 8.610 14.940 ;
        RECT 9.210 14.890 9.710 15.280 ;
        RECT 8.160 14.670 9.710 14.890 ;
        RECT 18.920 15.280 20.470 15.500 ;
        RECT 18.920 14.890 19.420 15.280 ;
        RECT 20.020 15.230 20.470 15.280 ;
        RECT 20.850 15.230 21.280 15.290 ;
        RECT 21.660 15.280 23.210 15.500 ;
        RECT 25.960 15.430 26.370 15.860 ;
        RECT 26.760 15.760 27.210 15.860 ;
        RECT 28.420 16.100 28.870 16.210 ;
        RECT 30.270 16.100 30.720 16.210 ;
        RECT 28.420 15.860 30.720 16.100 ;
        RECT 28.420 15.760 28.870 15.860 ;
        RECT 29.260 15.430 29.670 15.860 ;
        RECT 30.270 15.790 30.720 15.860 ;
        RECT 31.670 16.100 32.120 16.180 ;
        RECT 32.720 16.100 33.130 16.540 ;
        RECT 33.520 16.100 33.970 16.210 ;
        RECT 31.670 15.860 33.970 16.100 ;
        RECT 31.670 15.760 32.120 15.860 ;
        RECT 33.520 15.760 33.970 15.860 ;
        RECT 35.160 16.100 35.610 16.210 ;
        RECT 36.000 16.100 36.410 16.540 ;
        RECT 39.180 16.270 39.630 16.550 ;
        RECT 43.000 16.270 43.450 16.550 ;
        RECT 52.680 16.750 56.950 16.760 ;
        RECT 52.680 16.550 54.210 16.750 ;
        RECT 54.590 16.680 55.040 16.750 ;
        RECT 55.420 16.550 56.950 16.750 ;
        RECT 37.010 16.100 37.460 16.180 ;
        RECT 35.160 15.860 37.460 16.100 ;
        RECT 35.160 15.760 35.610 15.860 ;
        RECT 37.010 15.760 37.460 15.860 ;
        RECT 38.410 16.100 38.860 16.210 ;
        RECT 40.260 16.100 40.710 16.210 ;
        RECT 38.410 15.860 40.710 16.100 ;
        RECT 38.410 15.790 38.860 15.860 ;
        RECT 21.660 15.230 22.110 15.280 ;
        RECT 20.020 14.940 22.110 15.230 ;
        RECT 20.020 14.890 20.470 14.940 ;
        RECT 3.270 14.310 3.720 14.380 ;
        RECT 1.420 14.070 3.720 14.310 ;
        RECT 1.420 13.960 1.870 14.070 ;
        RECT 3.270 13.960 3.720 14.070 ;
        RECT 4.670 14.310 5.120 14.410 ;
        RECT 6.520 14.310 6.970 14.410 ;
        RECT 4.670 14.070 6.970 14.310 ;
        RECT 4.670 13.990 5.120 14.070 ;
        RECT 5.720 13.630 6.130 14.070 ;
        RECT 6.520 13.960 6.970 14.070 ;
        RECT 8.160 14.310 8.610 14.410 ;
        RECT 10.010 14.310 10.460 14.410 ;
        RECT 8.160 14.070 10.460 14.310 ;
        RECT 8.160 13.960 8.610 14.070 ;
        RECT 9.000 13.630 9.410 14.070 ;
        RECT 10.010 13.990 10.460 14.070 ;
        RECT 11.410 14.310 11.860 14.380 ;
        RECT 12.460 14.310 12.870 14.740 ;
        RECT 13.260 14.310 13.710 14.410 ;
        RECT 11.410 14.070 13.710 14.310 ;
        RECT 11.410 13.960 11.860 14.070 ;
        RECT 13.260 13.960 13.710 14.070 ;
        RECT 14.920 14.310 15.370 14.410 ;
        RECT 15.760 14.310 16.170 14.740 ;
        RECT 18.920 14.670 20.470 14.890 ;
        RECT 20.850 14.880 21.280 14.940 ;
        RECT 21.660 14.890 22.110 14.940 ;
        RECT 22.710 14.890 23.210 15.280 ;
        RECT 21.660 14.670 23.210 14.890 ;
        RECT 32.420 15.280 33.970 15.500 ;
        RECT 32.420 14.890 32.920 15.280 ;
        RECT 33.520 15.230 33.970 15.280 ;
        RECT 34.350 15.230 34.780 15.290 ;
        RECT 35.160 15.280 36.710 15.500 ;
        RECT 39.460 15.430 39.870 15.860 ;
        RECT 40.260 15.760 40.710 15.860 ;
        RECT 41.920 16.100 42.370 16.210 ;
        RECT 43.770 16.100 44.220 16.210 ;
        RECT 41.920 15.860 44.220 16.100 ;
        RECT 41.920 15.760 42.370 15.860 ;
        RECT 42.760 15.430 43.170 15.860 ;
        RECT 43.770 15.790 44.220 15.860 ;
        RECT 45.170 16.100 45.620 16.180 ;
        RECT 46.220 16.100 46.630 16.540 ;
        RECT 47.020 16.100 47.470 16.210 ;
        RECT 45.170 15.860 47.470 16.100 ;
        RECT 45.170 15.760 45.620 15.860 ;
        RECT 47.020 15.760 47.470 15.860 ;
        RECT 48.660 16.100 49.110 16.210 ;
        RECT 49.500 16.100 49.910 16.540 ;
        RECT 52.680 16.270 53.130 16.550 ;
        RECT 56.500 16.270 56.950 16.550 ;
        RECT 66.180 16.550 67.710 16.760 ;
        RECT 68.090 16.680 68.540 16.770 ;
        RECT 68.920 16.760 69.370 16.770 ;
        RECT 80.760 17.020 81.210 17.120 ;
        RECT 81.590 17.020 82.040 17.110 ;
        RECT 82.420 17.020 82.870 17.120 ;
        RECT 80.760 16.770 82.870 17.020 ;
        RECT 80.760 16.760 81.210 16.770 ;
        RECT 68.920 16.550 70.450 16.760 ;
        RECT 50.510 16.100 50.960 16.180 ;
        RECT 48.660 15.860 50.960 16.100 ;
        RECT 48.660 15.760 49.110 15.860 ;
        RECT 50.510 15.760 50.960 15.860 ;
        RECT 51.910 16.100 52.360 16.210 ;
        RECT 53.760 16.100 54.210 16.210 ;
        RECT 51.910 15.860 54.210 16.100 ;
        RECT 51.910 15.790 52.360 15.860 ;
        RECT 35.160 15.230 35.610 15.280 ;
        RECT 33.520 14.940 35.610 15.230 ;
        RECT 33.520 14.890 33.970 14.940 ;
        RECT 16.770 14.310 17.220 14.380 ;
        RECT 14.920 14.070 17.220 14.310 ;
        RECT 14.920 13.960 15.370 14.070 ;
        RECT 16.770 13.960 17.220 14.070 ;
        RECT 18.170 14.310 18.620 14.410 ;
        RECT 20.020 14.310 20.470 14.410 ;
        RECT 18.170 14.070 20.470 14.310 ;
        RECT 18.170 13.990 18.620 14.070 ;
        RECT 12.180 13.620 12.630 13.900 ;
        RECT 16.000 13.620 16.450 13.900 ;
        RECT 19.220 13.630 19.630 14.070 ;
        RECT 20.020 13.960 20.470 14.070 ;
        RECT 21.660 14.310 22.110 14.410 ;
        RECT 23.510 14.310 23.960 14.410 ;
        RECT 21.660 14.070 23.960 14.310 ;
        RECT 21.660 13.960 22.110 14.070 ;
        RECT 22.500 13.630 22.910 14.070 ;
        RECT 23.510 13.990 23.960 14.070 ;
        RECT 24.910 14.310 25.360 14.380 ;
        RECT 25.960 14.310 26.370 14.740 ;
        RECT 26.760 14.310 27.210 14.410 ;
        RECT 24.910 14.070 27.210 14.310 ;
        RECT 24.910 13.960 25.360 14.070 ;
        RECT 26.760 13.960 27.210 14.070 ;
        RECT 28.420 14.310 28.870 14.410 ;
        RECT 29.260 14.310 29.670 14.740 ;
        RECT 32.420 14.670 33.970 14.890 ;
        RECT 34.350 14.880 34.780 14.940 ;
        RECT 35.160 14.890 35.610 14.940 ;
        RECT 36.210 14.890 36.710 15.280 ;
        RECT 35.160 14.670 36.710 14.890 ;
        RECT 45.920 15.280 47.470 15.500 ;
        RECT 45.920 14.890 46.420 15.280 ;
        RECT 47.020 15.230 47.470 15.280 ;
        RECT 47.850 15.230 48.280 15.290 ;
        RECT 48.660 15.280 50.210 15.500 ;
        RECT 52.960 15.430 53.370 15.860 ;
        RECT 53.760 15.760 54.210 15.860 ;
        RECT 55.420 16.100 55.870 16.210 ;
        RECT 57.270 16.100 57.720 16.210 ;
        RECT 55.420 15.860 57.720 16.100 ;
        RECT 55.420 15.760 55.870 15.860 ;
        RECT 56.260 15.430 56.670 15.860 ;
        RECT 57.270 15.790 57.720 15.860 ;
        RECT 58.670 16.100 59.120 16.180 ;
        RECT 59.720 16.100 60.130 16.540 ;
        RECT 60.520 16.100 60.970 16.210 ;
        RECT 58.670 15.860 60.970 16.100 ;
        RECT 58.670 15.760 59.120 15.860 ;
        RECT 60.520 15.760 60.970 15.860 ;
        RECT 62.160 16.100 62.610 16.210 ;
        RECT 63.000 16.100 63.410 16.540 ;
        RECT 66.180 16.270 66.630 16.550 ;
        RECT 70.000 16.270 70.450 16.550 ;
        RECT 79.680 16.550 81.210 16.760 ;
        RECT 81.590 16.680 82.040 16.770 ;
        RECT 82.420 16.760 82.870 16.770 ;
        RECT 94.260 17.020 94.710 17.120 ;
        RECT 95.090 17.020 95.540 17.110 ;
        RECT 95.920 17.020 96.370 17.120 ;
        RECT 94.260 16.770 96.370 17.020 ;
        RECT 94.260 16.760 94.710 16.770 ;
        RECT 82.420 16.550 83.950 16.760 ;
        RECT 64.010 16.100 64.460 16.180 ;
        RECT 62.160 15.860 64.460 16.100 ;
        RECT 62.160 15.760 62.610 15.860 ;
        RECT 64.010 15.760 64.460 15.860 ;
        RECT 65.410 16.100 65.860 16.210 ;
        RECT 67.260 16.100 67.710 16.210 ;
        RECT 65.410 15.860 67.710 16.100 ;
        RECT 65.410 15.790 65.860 15.860 ;
        RECT 48.660 15.230 49.110 15.280 ;
        RECT 47.020 14.940 49.110 15.230 ;
        RECT 47.020 14.890 47.470 14.940 ;
        RECT 30.270 14.310 30.720 14.380 ;
        RECT 28.420 14.070 30.720 14.310 ;
        RECT 28.420 13.960 28.870 14.070 ;
        RECT 30.270 13.960 30.720 14.070 ;
        RECT 31.670 14.310 32.120 14.410 ;
        RECT 33.520 14.310 33.970 14.410 ;
        RECT 31.670 14.070 33.970 14.310 ;
        RECT 31.670 13.990 32.120 14.070 ;
        RECT 12.180 13.410 13.710 13.620 ;
        RECT 14.090 13.410 14.540 13.500 ;
        RECT 14.920 13.410 16.450 13.620 ;
        RECT 25.680 13.620 26.130 13.900 ;
        RECT 29.500 13.620 29.950 13.900 ;
        RECT 32.720 13.630 33.130 14.070 ;
        RECT 33.520 13.960 33.970 14.070 ;
        RECT 35.160 14.310 35.610 14.410 ;
        RECT 37.010 14.310 37.460 14.410 ;
        RECT 35.160 14.070 37.460 14.310 ;
        RECT 35.160 13.960 35.610 14.070 ;
        RECT 36.000 13.630 36.410 14.070 ;
        RECT 37.010 13.990 37.460 14.070 ;
        RECT 38.410 14.310 38.860 14.380 ;
        RECT 39.460 14.310 39.870 14.740 ;
        RECT 40.260 14.310 40.710 14.410 ;
        RECT 38.410 14.070 40.710 14.310 ;
        RECT 38.410 13.960 38.860 14.070 ;
        RECT 40.260 13.960 40.710 14.070 ;
        RECT 41.920 14.310 42.370 14.410 ;
        RECT 42.760 14.310 43.170 14.740 ;
        RECT 45.920 14.670 47.470 14.890 ;
        RECT 47.850 14.880 48.280 14.940 ;
        RECT 48.660 14.890 49.110 14.940 ;
        RECT 49.710 14.890 50.210 15.280 ;
        RECT 48.660 14.670 50.210 14.890 ;
        RECT 59.420 15.280 60.970 15.500 ;
        RECT 59.420 14.890 59.920 15.280 ;
        RECT 60.520 15.230 60.970 15.280 ;
        RECT 61.350 15.230 61.780 15.290 ;
        RECT 62.160 15.280 63.710 15.500 ;
        RECT 66.460 15.430 66.870 15.860 ;
        RECT 67.260 15.760 67.710 15.860 ;
        RECT 68.920 16.100 69.370 16.210 ;
        RECT 70.770 16.100 71.220 16.210 ;
        RECT 68.920 15.860 71.220 16.100 ;
        RECT 68.920 15.760 69.370 15.860 ;
        RECT 69.760 15.430 70.170 15.860 ;
        RECT 70.770 15.790 71.220 15.860 ;
        RECT 72.170 16.100 72.620 16.180 ;
        RECT 73.220 16.100 73.630 16.540 ;
        RECT 74.020 16.100 74.470 16.210 ;
        RECT 72.170 15.860 74.470 16.100 ;
        RECT 72.170 15.760 72.620 15.860 ;
        RECT 74.020 15.760 74.470 15.860 ;
        RECT 75.660 16.100 76.110 16.210 ;
        RECT 76.500 16.100 76.910 16.540 ;
        RECT 79.680 16.270 80.130 16.550 ;
        RECT 83.500 16.270 83.950 16.550 ;
        RECT 93.180 16.550 94.710 16.760 ;
        RECT 95.090 16.680 95.540 16.770 ;
        RECT 95.920 16.760 96.370 16.770 ;
        RECT 107.760 17.070 108.210 17.120 ;
        RECT 108.590 17.070 109.040 17.110 ;
        RECT 109.420 17.070 109.870 17.120 ;
        RECT 107.760 16.760 109.870 17.070 ;
        RECT 121.260 17.020 121.710 17.120 ;
        RECT 122.090 17.020 122.540 17.110 ;
        RECT 122.920 17.020 123.370 17.120 ;
        RECT 121.260 16.770 123.370 17.020 ;
        RECT 121.260 16.760 121.710 16.770 ;
        RECT 95.920 16.550 97.450 16.760 ;
        RECT 77.510 16.100 77.960 16.180 ;
        RECT 75.660 15.860 77.960 16.100 ;
        RECT 75.660 15.760 76.110 15.860 ;
        RECT 77.510 15.760 77.960 15.860 ;
        RECT 78.910 16.100 79.360 16.210 ;
        RECT 80.760 16.100 81.210 16.210 ;
        RECT 78.910 15.860 81.210 16.100 ;
        RECT 78.910 15.790 79.360 15.860 ;
        RECT 62.160 15.230 62.610 15.280 ;
        RECT 60.520 14.940 62.610 15.230 ;
        RECT 60.520 14.890 60.970 14.940 ;
        RECT 43.770 14.310 44.220 14.380 ;
        RECT 41.920 14.070 44.220 14.310 ;
        RECT 41.920 13.960 42.370 14.070 ;
        RECT 43.770 13.960 44.220 14.070 ;
        RECT 45.170 14.310 45.620 14.410 ;
        RECT 47.020 14.310 47.470 14.410 ;
        RECT 45.170 14.070 47.470 14.310 ;
        RECT 45.170 13.990 45.620 14.070 ;
        RECT 25.680 13.410 27.210 13.620 ;
        RECT 27.590 13.410 28.040 13.500 ;
        RECT 28.420 13.410 29.950 13.620 ;
        RECT 39.180 13.620 39.630 13.900 ;
        RECT 43.000 13.620 43.450 13.900 ;
        RECT 46.220 13.630 46.630 14.070 ;
        RECT 47.020 13.960 47.470 14.070 ;
        RECT 48.660 14.310 49.110 14.410 ;
        RECT 50.510 14.310 50.960 14.410 ;
        RECT 48.660 14.070 50.960 14.310 ;
        RECT 48.660 13.960 49.110 14.070 ;
        RECT 49.500 13.630 49.910 14.070 ;
        RECT 50.510 13.990 50.960 14.070 ;
        RECT 51.910 14.310 52.360 14.380 ;
        RECT 52.960 14.310 53.370 14.740 ;
        RECT 53.760 14.310 54.210 14.410 ;
        RECT 51.910 14.070 54.210 14.310 ;
        RECT 51.910 13.960 52.360 14.070 ;
        RECT 53.760 13.960 54.210 14.070 ;
        RECT 55.420 14.310 55.870 14.410 ;
        RECT 56.260 14.310 56.670 14.740 ;
        RECT 59.420 14.670 60.970 14.890 ;
        RECT 61.350 14.880 61.780 14.940 ;
        RECT 62.160 14.890 62.610 14.940 ;
        RECT 63.210 14.890 63.710 15.280 ;
        RECT 62.160 14.670 63.710 14.890 ;
        RECT 72.920 15.280 74.470 15.500 ;
        RECT 72.920 14.890 73.420 15.280 ;
        RECT 74.020 15.230 74.470 15.280 ;
        RECT 74.850 15.230 75.280 15.290 ;
        RECT 75.660 15.280 77.210 15.500 ;
        RECT 79.960 15.430 80.370 15.860 ;
        RECT 80.760 15.760 81.210 15.860 ;
        RECT 82.420 16.100 82.870 16.210 ;
        RECT 84.270 16.100 84.720 16.210 ;
        RECT 82.420 15.860 84.720 16.100 ;
        RECT 82.420 15.760 82.870 15.860 ;
        RECT 83.260 15.430 83.670 15.860 ;
        RECT 84.270 15.790 84.720 15.860 ;
        RECT 85.670 16.100 86.120 16.180 ;
        RECT 86.720 16.100 87.130 16.540 ;
        RECT 87.520 16.100 87.970 16.210 ;
        RECT 85.670 15.860 87.970 16.100 ;
        RECT 85.670 15.760 86.120 15.860 ;
        RECT 87.520 15.760 87.970 15.860 ;
        RECT 89.160 16.100 89.610 16.210 ;
        RECT 90.000 16.100 90.410 16.540 ;
        RECT 93.180 16.270 93.630 16.550 ;
        RECT 97.000 16.270 97.450 16.550 ;
        RECT 106.680 16.750 110.950 16.760 ;
        RECT 106.680 16.550 108.210 16.750 ;
        RECT 108.590 16.680 109.040 16.750 ;
        RECT 109.420 16.550 110.950 16.750 ;
        RECT 91.010 16.100 91.460 16.180 ;
        RECT 89.160 15.860 91.460 16.100 ;
        RECT 89.160 15.760 89.610 15.860 ;
        RECT 91.010 15.760 91.460 15.860 ;
        RECT 92.410 16.100 92.860 16.210 ;
        RECT 94.260 16.100 94.710 16.210 ;
        RECT 92.410 15.860 94.710 16.100 ;
        RECT 92.410 15.790 92.860 15.860 ;
        RECT 75.660 15.230 76.110 15.280 ;
        RECT 74.020 14.940 76.110 15.230 ;
        RECT 74.020 14.890 74.470 14.940 ;
        RECT 57.270 14.310 57.720 14.380 ;
        RECT 55.420 14.070 57.720 14.310 ;
        RECT 55.420 13.960 55.870 14.070 ;
        RECT 57.270 13.960 57.720 14.070 ;
        RECT 58.670 14.310 59.120 14.410 ;
        RECT 60.520 14.310 60.970 14.410 ;
        RECT 58.670 14.070 60.970 14.310 ;
        RECT 58.670 13.990 59.120 14.070 ;
        RECT 39.180 13.410 40.710 13.620 ;
        RECT 41.090 13.410 41.540 13.500 ;
        RECT 41.920 13.410 43.450 13.620 ;
        RECT 52.680 13.620 53.130 13.900 ;
        RECT 56.500 13.620 56.950 13.900 ;
        RECT 59.720 13.630 60.130 14.070 ;
        RECT 60.520 13.960 60.970 14.070 ;
        RECT 62.160 14.310 62.610 14.410 ;
        RECT 64.010 14.310 64.460 14.410 ;
        RECT 62.160 14.070 64.460 14.310 ;
        RECT 62.160 13.960 62.610 14.070 ;
        RECT 63.000 13.630 63.410 14.070 ;
        RECT 64.010 13.990 64.460 14.070 ;
        RECT 65.410 14.310 65.860 14.380 ;
        RECT 66.460 14.310 66.870 14.740 ;
        RECT 67.260 14.310 67.710 14.410 ;
        RECT 65.410 14.070 67.710 14.310 ;
        RECT 65.410 13.960 65.860 14.070 ;
        RECT 67.260 13.960 67.710 14.070 ;
        RECT 68.920 14.310 69.370 14.410 ;
        RECT 69.760 14.310 70.170 14.740 ;
        RECT 72.920 14.670 74.470 14.890 ;
        RECT 74.850 14.880 75.280 14.940 ;
        RECT 75.660 14.890 76.110 14.940 ;
        RECT 76.710 14.890 77.210 15.280 ;
        RECT 75.660 14.670 77.210 14.890 ;
        RECT 86.420 15.280 87.970 15.500 ;
        RECT 86.420 14.890 86.920 15.280 ;
        RECT 87.520 15.230 87.970 15.280 ;
        RECT 88.350 15.230 88.780 15.290 ;
        RECT 89.160 15.280 90.710 15.500 ;
        RECT 93.460 15.430 93.870 15.860 ;
        RECT 94.260 15.760 94.710 15.860 ;
        RECT 95.920 16.100 96.370 16.210 ;
        RECT 97.770 16.100 98.220 16.210 ;
        RECT 95.920 15.860 98.220 16.100 ;
        RECT 95.920 15.760 96.370 15.860 ;
        RECT 96.760 15.430 97.170 15.860 ;
        RECT 97.770 15.790 98.220 15.860 ;
        RECT 99.170 16.100 99.620 16.180 ;
        RECT 100.220 16.100 100.630 16.540 ;
        RECT 101.020 16.100 101.470 16.210 ;
        RECT 99.170 15.860 101.470 16.100 ;
        RECT 99.170 15.760 99.620 15.860 ;
        RECT 101.020 15.760 101.470 15.860 ;
        RECT 102.660 16.100 103.110 16.210 ;
        RECT 103.500 16.100 103.910 16.540 ;
        RECT 106.680 16.270 107.130 16.550 ;
        RECT 110.500 16.270 110.950 16.550 ;
        RECT 120.180 16.550 121.710 16.760 ;
        RECT 122.090 16.680 122.540 16.770 ;
        RECT 122.920 16.760 123.370 16.770 ;
        RECT 134.760 17.020 135.210 17.120 ;
        RECT 135.590 17.020 136.040 17.110 ;
        RECT 136.420 17.020 136.870 17.120 ;
        RECT 134.760 16.770 136.870 17.020 ;
        RECT 134.760 16.760 135.210 16.770 ;
        RECT 122.920 16.550 124.450 16.760 ;
        RECT 104.510 16.100 104.960 16.180 ;
        RECT 102.660 15.860 104.960 16.100 ;
        RECT 102.660 15.760 103.110 15.860 ;
        RECT 104.510 15.760 104.960 15.860 ;
        RECT 105.910 16.100 106.360 16.210 ;
        RECT 107.760 16.100 108.210 16.210 ;
        RECT 105.910 15.860 108.210 16.100 ;
        RECT 105.910 15.790 106.360 15.860 ;
        RECT 89.160 15.230 89.610 15.280 ;
        RECT 87.520 14.940 89.610 15.230 ;
        RECT 87.520 14.890 87.970 14.940 ;
        RECT 70.770 14.310 71.220 14.380 ;
        RECT 68.920 14.070 71.220 14.310 ;
        RECT 68.920 13.960 69.370 14.070 ;
        RECT 70.770 13.960 71.220 14.070 ;
        RECT 72.170 14.310 72.620 14.410 ;
        RECT 74.020 14.310 74.470 14.410 ;
        RECT 72.170 14.070 74.470 14.310 ;
        RECT 72.170 13.990 72.620 14.070 ;
        RECT 52.680 13.410 54.210 13.620 ;
        RECT 54.590 13.410 55.040 13.500 ;
        RECT 55.420 13.410 56.950 13.620 ;
        RECT 66.180 13.620 66.630 13.900 ;
        RECT 70.000 13.620 70.450 13.900 ;
        RECT 73.220 13.630 73.630 14.070 ;
        RECT 74.020 13.960 74.470 14.070 ;
        RECT 75.660 14.310 76.110 14.410 ;
        RECT 77.510 14.310 77.960 14.410 ;
        RECT 75.660 14.070 77.960 14.310 ;
        RECT 75.660 13.960 76.110 14.070 ;
        RECT 76.500 13.630 76.910 14.070 ;
        RECT 77.510 13.990 77.960 14.070 ;
        RECT 78.910 14.310 79.360 14.380 ;
        RECT 79.960 14.310 80.370 14.740 ;
        RECT 80.760 14.310 81.210 14.410 ;
        RECT 78.910 14.070 81.210 14.310 ;
        RECT 78.910 13.960 79.360 14.070 ;
        RECT 80.760 13.960 81.210 14.070 ;
        RECT 82.420 14.310 82.870 14.410 ;
        RECT 83.260 14.310 83.670 14.740 ;
        RECT 86.420 14.670 87.970 14.890 ;
        RECT 88.350 14.880 88.780 14.940 ;
        RECT 89.160 14.890 89.610 14.940 ;
        RECT 90.210 14.890 90.710 15.280 ;
        RECT 89.160 14.670 90.710 14.890 ;
        RECT 99.920 15.280 101.470 15.500 ;
        RECT 99.920 14.890 100.420 15.280 ;
        RECT 101.020 15.230 101.470 15.280 ;
        RECT 101.850 15.230 102.280 15.290 ;
        RECT 102.660 15.280 104.210 15.500 ;
        RECT 106.960 15.430 107.370 15.860 ;
        RECT 107.760 15.760 108.210 15.860 ;
        RECT 109.420 16.100 109.870 16.210 ;
        RECT 111.270 16.100 111.720 16.210 ;
        RECT 109.420 15.860 111.720 16.100 ;
        RECT 109.420 15.760 109.870 15.860 ;
        RECT 110.260 15.430 110.670 15.860 ;
        RECT 111.270 15.790 111.720 15.860 ;
        RECT 112.670 16.100 113.120 16.180 ;
        RECT 113.720 16.100 114.130 16.540 ;
        RECT 114.520 16.100 114.970 16.210 ;
        RECT 112.670 15.860 114.970 16.100 ;
        RECT 112.670 15.760 113.120 15.860 ;
        RECT 114.520 15.760 114.970 15.860 ;
        RECT 116.160 16.100 116.610 16.210 ;
        RECT 117.000 16.100 117.410 16.540 ;
        RECT 120.180 16.270 120.630 16.550 ;
        RECT 124.000 16.270 124.450 16.550 ;
        RECT 133.680 16.550 135.210 16.760 ;
        RECT 135.590 16.680 136.040 16.770 ;
        RECT 136.420 16.760 136.870 16.770 ;
        RECT 148.260 17.020 148.710 17.120 ;
        RECT 149.090 17.020 149.540 17.110 ;
        RECT 149.920 17.020 150.370 17.120 ;
        RECT 148.260 16.770 150.370 17.020 ;
        RECT 148.260 16.760 148.710 16.770 ;
        RECT 136.420 16.550 137.950 16.760 ;
        RECT 118.010 16.100 118.460 16.180 ;
        RECT 116.160 15.860 118.460 16.100 ;
        RECT 116.160 15.760 116.610 15.860 ;
        RECT 118.010 15.760 118.460 15.860 ;
        RECT 119.410 16.100 119.860 16.210 ;
        RECT 121.260 16.100 121.710 16.210 ;
        RECT 119.410 15.860 121.710 16.100 ;
        RECT 119.410 15.790 119.860 15.860 ;
        RECT 102.660 15.230 103.110 15.280 ;
        RECT 101.020 14.940 103.110 15.230 ;
        RECT 101.020 14.890 101.470 14.940 ;
        RECT 84.270 14.310 84.720 14.380 ;
        RECT 82.420 14.070 84.720 14.310 ;
        RECT 82.420 13.960 82.870 14.070 ;
        RECT 84.270 13.960 84.720 14.070 ;
        RECT 85.670 14.310 86.120 14.410 ;
        RECT 87.520 14.310 87.970 14.410 ;
        RECT 85.670 14.070 87.970 14.310 ;
        RECT 85.670 13.990 86.120 14.070 ;
        RECT 66.180 13.410 67.710 13.620 ;
        RECT 68.090 13.410 68.540 13.500 ;
        RECT 68.920 13.410 70.450 13.620 ;
        RECT 79.680 13.620 80.130 13.900 ;
        RECT 83.500 13.620 83.950 13.900 ;
        RECT 86.720 13.630 87.130 14.070 ;
        RECT 87.520 13.960 87.970 14.070 ;
        RECT 89.160 14.310 89.610 14.410 ;
        RECT 91.010 14.310 91.460 14.410 ;
        RECT 89.160 14.070 91.460 14.310 ;
        RECT 89.160 13.960 89.610 14.070 ;
        RECT 90.000 13.630 90.410 14.070 ;
        RECT 91.010 13.990 91.460 14.070 ;
        RECT 92.410 14.310 92.860 14.380 ;
        RECT 93.460 14.310 93.870 14.740 ;
        RECT 94.260 14.310 94.710 14.410 ;
        RECT 92.410 14.070 94.710 14.310 ;
        RECT 92.410 13.960 92.860 14.070 ;
        RECT 94.260 13.960 94.710 14.070 ;
        RECT 95.920 14.310 96.370 14.410 ;
        RECT 96.760 14.310 97.170 14.740 ;
        RECT 99.920 14.670 101.470 14.890 ;
        RECT 101.850 14.880 102.280 14.940 ;
        RECT 102.660 14.890 103.110 14.940 ;
        RECT 103.710 14.890 104.210 15.280 ;
        RECT 102.660 14.670 104.210 14.890 ;
        RECT 113.420 15.280 114.970 15.500 ;
        RECT 113.420 14.890 113.920 15.280 ;
        RECT 114.520 15.230 114.970 15.280 ;
        RECT 115.350 15.230 115.780 15.290 ;
        RECT 116.160 15.280 117.710 15.500 ;
        RECT 120.460 15.430 120.870 15.860 ;
        RECT 121.260 15.760 121.710 15.860 ;
        RECT 122.920 16.100 123.370 16.210 ;
        RECT 124.770 16.100 125.220 16.210 ;
        RECT 122.920 15.860 125.220 16.100 ;
        RECT 122.920 15.760 123.370 15.860 ;
        RECT 123.760 15.430 124.170 15.860 ;
        RECT 124.770 15.790 125.220 15.860 ;
        RECT 126.170 16.100 126.620 16.180 ;
        RECT 127.220 16.100 127.630 16.540 ;
        RECT 128.020 16.100 128.470 16.210 ;
        RECT 126.170 15.860 128.470 16.100 ;
        RECT 126.170 15.760 126.620 15.860 ;
        RECT 128.020 15.760 128.470 15.860 ;
        RECT 129.660 16.100 130.110 16.210 ;
        RECT 130.500 16.100 130.910 16.540 ;
        RECT 133.680 16.270 134.130 16.550 ;
        RECT 137.500 16.270 137.950 16.550 ;
        RECT 147.180 16.550 148.710 16.760 ;
        RECT 149.090 16.680 149.540 16.770 ;
        RECT 149.920 16.760 150.370 16.770 ;
        RECT 161.760 17.070 162.210 17.120 ;
        RECT 162.590 17.070 163.040 17.110 ;
        RECT 163.420 17.070 163.870 17.120 ;
        RECT 161.760 16.760 163.870 17.070 ;
        RECT 175.260 17.020 175.710 17.120 ;
        RECT 176.090 17.020 176.540 17.110 ;
        RECT 176.920 17.020 177.370 17.120 ;
        RECT 175.260 16.770 177.370 17.020 ;
        RECT 175.260 16.760 175.710 16.770 ;
        RECT 149.920 16.550 151.450 16.760 ;
        RECT 131.510 16.100 131.960 16.180 ;
        RECT 129.660 15.860 131.960 16.100 ;
        RECT 129.660 15.760 130.110 15.860 ;
        RECT 131.510 15.760 131.960 15.860 ;
        RECT 132.910 16.100 133.360 16.210 ;
        RECT 134.760 16.100 135.210 16.210 ;
        RECT 132.910 15.860 135.210 16.100 ;
        RECT 132.910 15.790 133.360 15.860 ;
        RECT 116.160 15.230 116.610 15.280 ;
        RECT 114.520 14.940 116.610 15.230 ;
        RECT 114.520 14.890 114.970 14.940 ;
        RECT 97.770 14.310 98.220 14.380 ;
        RECT 95.920 14.070 98.220 14.310 ;
        RECT 95.920 13.960 96.370 14.070 ;
        RECT 97.770 13.960 98.220 14.070 ;
        RECT 99.170 14.310 99.620 14.410 ;
        RECT 101.020 14.310 101.470 14.410 ;
        RECT 99.170 14.070 101.470 14.310 ;
        RECT 99.170 13.990 99.620 14.070 ;
        RECT 79.680 13.410 81.210 13.620 ;
        RECT 81.590 13.410 82.040 13.500 ;
        RECT 82.420 13.410 83.950 13.620 ;
        RECT 93.180 13.620 93.630 13.900 ;
        RECT 97.000 13.620 97.450 13.900 ;
        RECT 100.220 13.630 100.630 14.070 ;
        RECT 101.020 13.960 101.470 14.070 ;
        RECT 102.660 14.310 103.110 14.410 ;
        RECT 104.510 14.310 104.960 14.410 ;
        RECT 102.660 14.070 104.960 14.310 ;
        RECT 102.660 13.960 103.110 14.070 ;
        RECT 103.500 13.630 103.910 14.070 ;
        RECT 104.510 13.990 104.960 14.070 ;
        RECT 105.910 14.310 106.360 14.380 ;
        RECT 106.960 14.310 107.370 14.740 ;
        RECT 107.760 14.310 108.210 14.410 ;
        RECT 105.910 14.070 108.210 14.310 ;
        RECT 105.910 13.960 106.360 14.070 ;
        RECT 107.760 13.960 108.210 14.070 ;
        RECT 109.420 14.310 109.870 14.410 ;
        RECT 110.260 14.310 110.670 14.740 ;
        RECT 113.420 14.670 114.970 14.890 ;
        RECT 115.350 14.880 115.780 14.940 ;
        RECT 116.160 14.890 116.610 14.940 ;
        RECT 117.210 14.890 117.710 15.280 ;
        RECT 116.160 14.670 117.710 14.890 ;
        RECT 126.920 15.280 128.470 15.500 ;
        RECT 126.920 14.890 127.420 15.280 ;
        RECT 128.020 15.230 128.470 15.280 ;
        RECT 128.850 15.230 129.280 15.290 ;
        RECT 129.660 15.280 131.210 15.500 ;
        RECT 133.960 15.430 134.370 15.860 ;
        RECT 134.760 15.760 135.210 15.860 ;
        RECT 136.420 16.100 136.870 16.210 ;
        RECT 138.270 16.100 138.720 16.210 ;
        RECT 136.420 15.860 138.720 16.100 ;
        RECT 136.420 15.760 136.870 15.860 ;
        RECT 137.260 15.430 137.670 15.860 ;
        RECT 138.270 15.790 138.720 15.860 ;
        RECT 139.670 16.100 140.120 16.180 ;
        RECT 140.720 16.100 141.130 16.540 ;
        RECT 141.520 16.100 141.970 16.210 ;
        RECT 139.670 15.860 141.970 16.100 ;
        RECT 139.670 15.760 140.120 15.860 ;
        RECT 141.520 15.760 141.970 15.860 ;
        RECT 143.160 16.100 143.610 16.210 ;
        RECT 144.000 16.100 144.410 16.540 ;
        RECT 147.180 16.270 147.630 16.550 ;
        RECT 151.000 16.270 151.450 16.550 ;
        RECT 160.680 16.750 164.950 16.760 ;
        RECT 160.680 16.550 162.210 16.750 ;
        RECT 162.590 16.680 163.040 16.750 ;
        RECT 163.420 16.550 164.950 16.750 ;
        RECT 145.010 16.100 145.460 16.180 ;
        RECT 143.160 15.860 145.460 16.100 ;
        RECT 143.160 15.760 143.610 15.860 ;
        RECT 145.010 15.760 145.460 15.860 ;
        RECT 146.410 16.100 146.860 16.210 ;
        RECT 148.260 16.100 148.710 16.210 ;
        RECT 146.410 15.860 148.710 16.100 ;
        RECT 146.410 15.790 146.860 15.860 ;
        RECT 129.660 15.230 130.110 15.280 ;
        RECT 128.020 14.940 130.110 15.230 ;
        RECT 128.020 14.890 128.470 14.940 ;
        RECT 111.270 14.310 111.720 14.380 ;
        RECT 109.420 14.070 111.720 14.310 ;
        RECT 109.420 13.960 109.870 14.070 ;
        RECT 111.270 13.960 111.720 14.070 ;
        RECT 112.670 14.310 113.120 14.410 ;
        RECT 114.520 14.310 114.970 14.410 ;
        RECT 112.670 14.070 114.970 14.310 ;
        RECT 112.670 13.990 113.120 14.070 ;
        RECT 93.180 13.410 94.710 13.620 ;
        RECT 95.090 13.410 95.540 13.500 ;
        RECT 95.920 13.410 97.450 13.620 ;
        RECT 106.680 13.620 107.130 13.900 ;
        RECT 110.500 13.620 110.950 13.900 ;
        RECT 113.720 13.630 114.130 14.070 ;
        RECT 114.520 13.960 114.970 14.070 ;
        RECT 116.160 14.310 116.610 14.410 ;
        RECT 118.010 14.310 118.460 14.410 ;
        RECT 116.160 14.070 118.460 14.310 ;
        RECT 116.160 13.960 116.610 14.070 ;
        RECT 117.000 13.630 117.410 14.070 ;
        RECT 118.010 13.990 118.460 14.070 ;
        RECT 119.410 14.310 119.860 14.380 ;
        RECT 120.460 14.310 120.870 14.740 ;
        RECT 121.260 14.310 121.710 14.410 ;
        RECT 119.410 14.070 121.710 14.310 ;
        RECT 119.410 13.960 119.860 14.070 ;
        RECT 121.260 13.960 121.710 14.070 ;
        RECT 122.920 14.310 123.370 14.410 ;
        RECT 123.760 14.310 124.170 14.740 ;
        RECT 126.920 14.670 128.470 14.890 ;
        RECT 128.850 14.880 129.280 14.940 ;
        RECT 129.660 14.890 130.110 14.940 ;
        RECT 130.710 14.890 131.210 15.280 ;
        RECT 129.660 14.670 131.210 14.890 ;
        RECT 140.420 15.280 141.970 15.500 ;
        RECT 140.420 14.890 140.920 15.280 ;
        RECT 141.520 15.230 141.970 15.280 ;
        RECT 142.350 15.230 142.780 15.290 ;
        RECT 143.160 15.280 144.710 15.500 ;
        RECT 147.460 15.430 147.870 15.860 ;
        RECT 148.260 15.760 148.710 15.860 ;
        RECT 149.920 16.100 150.370 16.210 ;
        RECT 151.770 16.100 152.220 16.210 ;
        RECT 149.920 15.860 152.220 16.100 ;
        RECT 149.920 15.760 150.370 15.860 ;
        RECT 150.760 15.430 151.170 15.860 ;
        RECT 151.770 15.790 152.220 15.860 ;
        RECT 153.170 16.100 153.620 16.180 ;
        RECT 154.220 16.100 154.630 16.540 ;
        RECT 155.020 16.100 155.470 16.210 ;
        RECT 153.170 15.860 155.470 16.100 ;
        RECT 153.170 15.760 153.620 15.860 ;
        RECT 155.020 15.760 155.470 15.860 ;
        RECT 156.660 16.100 157.110 16.210 ;
        RECT 157.500 16.100 157.910 16.540 ;
        RECT 160.680 16.270 161.130 16.550 ;
        RECT 164.500 16.270 164.950 16.550 ;
        RECT 174.180 16.550 175.710 16.760 ;
        RECT 176.090 16.680 176.540 16.770 ;
        RECT 176.920 16.760 177.370 16.770 ;
        RECT 188.760 17.020 189.210 17.120 ;
        RECT 189.590 17.020 190.040 17.110 ;
        RECT 190.420 17.020 190.870 17.120 ;
        RECT 188.760 16.770 190.870 17.020 ;
        RECT 188.760 16.760 189.210 16.770 ;
        RECT 176.920 16.550 178.450 16.760 ;
        RECT 158.510 16.100 158.960 16.180 ;
        RECT 156.660 15.860 158.960 16.100 ;
        RECT 156.660 15.760 157.110 15.860 ;
        RECT 158.510 15.760 158.960 15.860 ;
        RECT 159.910 16.100 160.360 16.210 ;
        RECT 161.760 16.100 162.210 16.210 ;
        RECT 159.910 15.860 162.210 16.100 ;
        RECT 159.910 15.790 160.360 15.860 ;
        RECT 143.160 15.230 143.610 15.280 ;
        RECT 141.520 14.940 143.610 15.230 ;
        RECT 141.520 14.890 141.970 14.940 ;
        RECT 124.770 14.310 125.220 14.380 ;
        RECT 122.920 14.070 125.220 14.310 ;
        RECT 122.920 13.960 123.370 14.070 ;
        RECT 124.770 13.960 125.220 14.070 ;
        RECT 126.170 14.310 126.620 14.410 ;
        RECT 128.020 14.310 128.470 14.410 ;
        RECT 126.170 14.070 128.470 14.310 ;
        RECT 126.170 13.990 126.620 14.070 ;
        RECT 106.680 13.410 108.210 13.620 ;
        RECT 108.590 13.410 109.040 13.500 ;
        RECT 109.420 13.410 110.950 13.620 ;
        RECT 120.180 13.620 120.630 13.900 ;
        RECT 124.000 13.620 124.450 13.900 ;
        RECT 127.220 13.630 127.630 14.070 ;
        RECT 128.020 13.960 128.470 14.070 ;
        RECT 129.660 14.310 130.110 14.410 ;
        RECT 131.510 14.310 131.960 14.410 ;
        RECT 129.660 14.070 131.960 14.310 ;
        RECT 129.660 13.960 130.110 14.070 ;
        RECT 130.500 13.630 130.910 14.070 ;
        RECT 131.510 13.990 131.960 14.070 ;
        RECT 132.910 14.310 133.360 14.380 ;
        RECT 133.960 14.310 134.370 14.740 ;
        RECT 134.760 14.310 135.210 14.410 ;
        RECT 132.910 14.070 135.210 14.310 ;
        RECT 132.910 13.960 133.360 14.070 ;
        RECT 134.760 13.960 135.210 14.070 ;
        RECT 136.420 14.310 136.870 14.410 ;
        RECT 137.260 14.310 137.670 14.740 ;
        RECT 140.420 14.670 141.970 14.890 ;
        RECT 142.350 14.880 142.780 14.940 ;
        RECT 143.160 14.890 143.610 14.940 ;
        RECT 144.210 14.890 144.710 15.280 ;
        RECT 143.160 14.670 144.710 14.890 ;
        RECT 153.920 15.280 155.470 15.500 ;
        RECT 153.920 14.890 154.420 15.280 ;
        RECT 155.020 15.230 155.470 15.280 ;
        RECT 155.850 15.230 156.280 15.290 ;
        RECT 156.660 15.280 158.210 15.500 ;
        RECT 160.960 15.430 161.370 15.860 ;
        RECT 161.760 15.760 162.210 15.860 ;
        RECT 163.420 16.100 163.870 16.210 ;
        RECT 165.270 16.100 165.720 16.210 ;
        RECT 163.420 15.860 165.720 16.100 ;
        RECT 163.420 15.760 163.870 15.860 ;
        RECT 164.260 15.430 164.670 15.860 ;
        RECT 165.270 15.790 165.720 15.860 ;
        RECT 166.670 16.100 167.120 16.180 ;
        RECT 167.720 16.100 168.130 16.540 ;
        RECT 168.520 16.100 168.970 16.210 ;
        RECT 166.670 15.860 168.970 16.100 ;
        RECT 166.670 15.760 167.120 15.860 ;
        RECT 168.520 15.760 168.970 15.860 ;
        RECT 170.160 16.100 170.610 16.210 ;
        RECT 171.000 16.100 171.410 16.540 ;
        RECT 174.180 16.270 174.630 16.550 ;
        RECT 178.000 16.270 178.450 16.550 ;
        RECT 187.680 16.550 189.210 16.760 ;
        RECT 189.590 16.680 190.040 16.770 ;
        RECT 190.420 16.760 190.870 16.770 ;
        RECT 202.260 17.020 202.710 17.120 ;
        RECT 203.090 17.020 203.540 17.110 ;
        RECT 203.920 17.020 204.370 17.120 ;
        RECT 202.260 16.770 204.370 17.020 ;
        RECT 202.260 16.760 202.710 16.770 ;
        RECT 190.420 16.550 191.950 16.760 ;
        RECT 172.010 16.100 172.460 16.180 ;
        RECT 170.160 15.860 172.460 16.100 ;
        RECT 170.160 15.760 170.610 15.860 ;
        RECT 172.010 15.760 172.460 15.860 ;
        RECT 173.410 16.100 173.860 16.210 ;
        RECT 175.260 16.100 175.710 16.210 ;
        RECT 173.410 15.860 175.710 16.100 ;
        RECT 173.410 15.790 173.860 15.860 ;
        RECT 156.660 15.230 157.110 15.280 ;
        RECT 155.020 14.940 157.110 15.230 ;
        RECT 155.020 14.890 155.470 14.940 ;
        RECT 138.270 14.310 138.720 14.380 ;
        RECT 136.420 14.070 138.720 14.310 ;
        RECT 136.420 13.960 136.870 14.070 ;
        RECT 138.270 13.960 138.720 14.070 ;
        RECT 139.670 14.310 140.120 14.410 ;
        RECT 141.520 14.310 141.970 14.410 ;
        RECT 139.670 14.070 141.970 14.310 ;
        RECT 139.670 13.990 140.120 14.070 ;
        RECT 120.180 13.410 121.710 13.620 ;
        RECT 122.090 13.410 122.540 13.500 ;
        RECT 122.920 13.410 124.450 13.620 ;
        RECT 133.680 13.620 134.130 13.900 ;
        RECT 137.500 13.620 137.950 13.900 ;
        RECT 140.720 13.630 141.130 14.070 ;
        RECT 141.520 13.960 141.970 14.070 ;
        RECT 143.160 14.310 143.610 14.410 ;
        RECT 145.010 14.310 145.460 14.410 ;
        RECT 143.160 14.070 145.460 14.310 ;
        RECT 143.160 13.960 143.610 14.070 ;
        RECT 144.000 13.630 144.410 14.070 ;
        RECT 145.010 13.990 145.460 14.070 ;
        RECT 146.410 14.310 146.860 14.380 ;
        RECT 147.460 14.310 147.870 14.740 ;
        RECT 148.260 14.310 148.710 14.410 ;
        RECT 146.410 14.070 148.710 14.310 ;
        RECT 146.410 13.960 146.860 14.070 ;
        RECT 148.260 13.960 148.710 14.070 ;
        RECT 149.920 14.310 150.370 14.410 ;
        RECT 150.760 14.310 151.170 14.740 ;
        RECT 153.920 14.670 155.470 14.890 ;
        RECT 155.850 14.880 156.280 14.940 ;
        RECT 156.660 14.890 157.110 14.940 ;
        RECT 157.710 14.890 158.210 15.280 ;
        RECT 156.660 14.670 158.210 14.890 ;
        RECT 167.420 15.280 168.970 15.500 ;
        RECT 167.420 14.890 167.920 15.280 ;
        RECT 168.520 15.230 168.970 15.280 ;
        RECT 169.350 15.230 169.780 15.290 ;
        RECT 170.160 15.280 171.710 15.500 ;
        RECT 174.460 15.430 174.870 15.860 ;
        RECT 175.260 15.760 175.710 15.860 ;
        RECT 176.920 16.100 177.370 16.210 ;
        RECT 178.770 16.100 179.220 16.210 ;
        RECT 176.920 15.860 179.220 16.100 ;
        RECT 176.920 15.760 177.370 15.860 ;
        RECT 177.760 15.430 178.170 15.860 ;
        RECT 178.770 15.790 179.220 15.860 ;
        RECT 180.170 16.100 180.620 16.180 ;
        RECT 181.220 16.100 181.630 16.540 ;
        RECT 182.020 16.100 182.470 16.210 ;
        RECT 180.170 15.860 182.470 16.100 ;
        RECT 180.170 15.760 180.620 15.860 ;
        RECT 182.020 15.760 182.470 15.860 ;
        RECT 183.660 16.100 184.110 16.210 ;
        RECT 184.500 16.100 184.910 16.540 ;
        RECT 187.680 16.270 188.130 16.550 ;
        RECT 191.500 16.270 191.950 16.550 ;
        RECT 201.180 16.550 202.710 16.760 ;
        RECT 203.090 16.680 203.540 16.770 ;
        RECT 203.920 16.760 204.370 16.770 ;
        RECT 215.760 17.020 216.210 17.120 ;
        RECT 216.590 17.070 217.030 17.110 ;
        RECT 216.590 17.020 217.690 17.070 ;
        RECT 215.760 16.770 217.690 17.020 ;
        RECT 215.760 16.760 216.210 16.770 ;
        RECT 203.920 16.550 205.450 16.760 ;
        RECT 185.510 16.100 185.960 16.180 ;
        RECT 183.660 15.860 185.960 16.100 ;
        RECT 183.660 15.760 184.110 15.860 ;
        RECT 185.510 15.760 185.960 15.860 ;
        RECT 186.910 16.100 187.360 16.210 ;
        RECT 188.760 16.100 189.210 16.210 ;
        RECT 186.910 15.860 189.210 16.100 ;
        RECT 186.910 15.790 187.360 15.860 ;
        RECT 170.160 15.230 170.610 15.280 ;
        RECT 168.520 14.940 170.610 15.230 ;
        RECT 168.520 14.890 168.970 14.940 ;
        RECT 151.770 14.310 152.220 14.380 ;
        RECT 149.920 14.070 152.220 14.310 ;
        RECT 149.920 13.960 150.370 14.070 ;
        RECT 151.770 13.960 152.220 14.070 ;
        RECT 153.170 14.310 153.620 14.410 ;
        RECT 155.020 14.310 155.470 14.410 ;
        RECT 153.170 14.070 155.470 14.310 ;
        RECT 153.170 13.990 153.620 14.070 ;
        RECT 133.680 13.410 135.210 13.620 ;
        RECT 135.590 13.410 136.040 13.500 ;
        RECT 136.420 13.410 137.950 13.620 ;
        RECT 147.180 13.620 147.630 13.900 ;
        RECT 151.000 13.620 151.450 13.900 ;
        RECT 154.220 13.630 154.630 14.070 ;
        RECT 155.020 13.960 155.470 14.070 ;
        RECT 156.660 14.310 157.110 14.410 ;
        RECT 158.510 14.310 158.960 14.410 ;
        RECT 156.660 14.070 158.960 14.310 ;
        RECT 156.660 13.960 157.110 14.070 ;
        RECT 157.500 13.630 157.910 14.070 ;
        RECT 158.510 13.990 158.960 14.070 ;
        RECT 159.910 14.310 160.360 14.380 ;
        RECT 160.960 14.310 161.370 14.740 ;
        RECT 161.760 14.310 162.210 14.410 ;
        RECT 159.910 14.070 162.210 14.310 ;
        RECT 159.910 13.960 160.360 14.070 ;
        RECT 161.760 13.960 162.210 14.070 ;
        RECT 163.420 14.310 163.870 14.410 ;
        RECT 164.260 14.310 164.670 14.740 ;
        RECT 167.420 14.670 168.970 14.890 ;
        RECT 169.350 14.880 169.780 14.940 ;
        RECT 170.160 14.890 170.610 14.940 ;
        RECT 171.210 14.890 171.710 15.280 ;
        RECT 170.160 14.670 171.710 14.890 ;
        RECT 180.920 15.280 182.470 15.500 ;
        RECT 180.920 14.890 181.420 15.280 ;
        RECT 182.020 15.230 182.470 15.280 ;
        RECT 182.850 15.230 183.280 15.290 ;
        RECT 183.660 15.280 185.210 15.500 ;
        RECT 187.960 15.430 188.370 15.860 ;
        RECT 188.760 15.760 189.210 15.860 ;
        RECT 190.420 16.100 190.870 16.210 ;
        RECT 192.270 16.100 192.720 16.210 ;
        RECT 190.420 15.860 192.720 16.100 ;
        RECT 190.420 15.760 190.870 15.860 ;
        RECT 191.260 15.430 191.670 15.860 ;
        RECT 192.270 15.790 192.720 15.860 ;
        RECT 193.670 16.100 194.120 16.180 ;
        RECT 194.720 16.100 195.130 16.540 ;
        RECT 195.520 16.100 195.970 16.210 ;
        RECT 193.670 15.860 195.970 16.100 ;
        RECT 193.670 15.760 194.120 15.860 ;
        RECT 195.520 15.760 195.970 15.860 ;
        RECT 197.160 16.100 197.610 16.210 ;
        RECT 198.000 16.100 198.410 16.540 ;
        RECT 201.180 16.270 201.630 16.550 ;
        RECT 205.000 16.270 205.450 16.550 ;
        RECT 214.680 16.550 216.210 16.760 ;
        RECT 216.590 16.750 217.690 16.770 ;
        RECT 216.590 16.680 217.030 16.750 ;
        RECT 199.010 16.100 199.460 16.180 ;
        RECT 197.160 15.860 199.460 16.100 ;
        RECT 197.160 15.760 197.610 15.860 ;
        RECT 199.010 15.760 199.460 15.860 ;
        RECT 200.410 16.100 200.860 16.210 ;
        RECT 202.260 16.100 202.710 16.210 ;
        RECT 200.410 15.860 202.710 16.100 ;
        RECT 200.410 15.790 200.860 15.860 ;
        RECT 183.660 15.230 184.110 15.280 ;
        RECT 182.020 14.940 184.110 15.230 ;
        RECT 182.020 14.890 182.470 14.940 ;
        RECT 165.270 14.310 165.720 14.380 ;
        RECT 163.420 14.070 165.720 14.310 ;
        RECT 163.420 13.960 163.870 14.070 ;
        RECT 165.270 13.960 165.720 14.070 ;
        RECT 166.670 14.310 167.120 14.410 ;
        RECT 168.520 14.310 168.970 14.410 ;
        RECT 166.670 14.070 168.970 14.310 ;
        RECT 166.670 13.990 167.120 14.070 ;
        RECT 147.180 13.410 148.710 13.620 ;
        RECT 149.090 13.410 149.540 13.500 ;
        RECT 149.920 13.410 151.450 13.620 ;
        RECT 160.680 13.620 161.130 13.900 ;
        RECT 164.500 13.620 164.950 13.900 ;
        RECT 167.720 13.630 168.130 14.070 ;
        RECT 168.520 13.960 168.970 14.070 ;
        RECT 170.160 14.310 170.610 14.410 ;
        RECT 172.010 14.310 172.460 14.410 ;
        RECT 170.160 14.070 172.460 14.310 ;
        RECT 170.160 13.960 170.610 14.070 ;
        RECT 171.000 13.630 171.410 14.070 ;
        RECT 172.010 13.990 172.460 14.070 ;
        RECT 173.410 14.310 173.860 14.380 ;
        RECT 174.460 14.310 174.870 14.740 ;
        RECT 175.260 14.310 175.710 14.410 ;
        RECT 173.410 14.070 175.710 14.310 ;
        RECT 173.410 13.960 173.860 14.070 ;
        RECT 175.260 13.960 175.710 14.070 ;
        RECT 176.920 14.310 177.370 14.410 ;
        RECT 177.760 14.310 178.170 14.740 ;
        RECT 180.920 14.670 182.470 14.890 ;
        RECT 182.850 14.880 183.280 14.940 ;
        RECT 183.660 14.890 184.110 14.940 ;
        RECT 184.710 14.890 185.210 15.280 ;
        RECT 183.660 14.670 185.210 14.890 ;
        RECT 194.420 15.280 195.970 15.500 ;
        RECT 194.420 14.890 194.920 15.280 ;
        RECT 195.520 15.230 195.970 15.280 ;
        RECT 196.350 15.230 196.780 15.290 ;
        RECT 197.160 15.280 198.710 15.500 ;
        RECT 201.460 15.430 201.870 15.860 ;
        RECT 202.260 15.760 202.710 15.860 ;
        RECT 203.920 16.100 204.370 16.210 ;
        RECT 205.770 16.100 206.220 16.210 ;
        RECT 203.920 15.860 206.220 16.100 ;
        RECT 203.920 15.760 204.370 15.860 ;
        RECT 204.760 15.430 205.170 15.860 ;
        RECT 205.770 15.790 206.220 15.860 ;
        RECT 207.170 16.100 207.620 16.180 ;
        RECT 208.220 16.100 208.630 16.540 ;
        RECT 209.020 16.100 209.470 16.210 ;
        RECT 207.170 15.860 209.470 16.100 ;
        RECT 207.170 15.760 207.620 15.860 ;
        RECT 209.020 15.760 209.470 15.860 ;
        RECT 210.660 16.100 211.110 16.210 ;
        RECT 211.500 16.100 211.910 16.540 ;
        RECT 214.680 16.270 215.130 16.550 ;
        RECT 212.510 16.100 212.960 16.180 ;
        RECT 210.660 15.860 212.960 16.100 ;
        RECT 210.660 15.760 211.110 15.860 ;
        RECT 212.510 15.760 212.960 15.860 ;
        RECT 213.910 16.100 214.360 16.210 ;
        RECT 215.760 16.100 216.210 16.210 ;
        RECT 213.910 15.860 216.210 16.100 ;
        RECT 213.910 15.790 214.360 15.860 ;
        RECT 197.160 15.230 197.610 15.280 ;
        RECT 195.520 14.940 197.610 15.230 ;
        RECT 195.520 14.890 195.970 14.940 ;
        RECT 178.770 14.310 179.220 14.380 ;
        RECT 176.920 14.070 179.220 14.310 ;
        RECT 176.920 13.960 177.370 14.070 ;
        RECT 178.770 13.960 179.220 14.070 ;
        RECT 180.170 14.310 180.620 14.410 ;
        RECT 182.020 14.310 182.470 14.410 ;
        RECT 180.170 14.070 182.470 14.310 ;
        RECT 180.170 13.990 180.620 14.070 ;
        RECT 160.680 13.410 162.210 13.620 ;
        RECT 162.590 13.410 163.040 13.500 ;
        RECT 163.420 13.410 164.950 13.620 ;
        RECT 174.180 13.620 174.630 13.900 ;
        RECT 178.000 13.620 178.450 13.900 ;
        RECT 181.220 13.630 181.630 14.070 ;
        RECT 182.020 13.960 182.470 14.070 ;
        RECT 183.660 14.310 184.110 14.410 ;
        RECT 185.510 14.310 185.960 14.410 ;
        RECT 183.660 14.070 185.960 14.310 ;
        RECT 183.660 13.960 184.110 14.070 ;
        RECT 184.500 13.630 184.910 14.070 ;
        RECT 185.510 13.990 185.960 14.070 ;
        RECT 186.910 14.310 187.360 14.380 ;
        RECT 187.960 14.310 188.370 14.740 ;
        RECT 188.760 14.310 189.210 14.410 ;
        RECT 186.910 14.070 189.210 14.310 ;
        RECT 186.910 13.960 187.360 14.070 ;
        RECT 188.760 13.960 189.210 14.070 ;
        RECT 190.420 14.310 190.870 14.410 ;
        RECT 191.260 14.310 191.670 14.740 ;
        RECT 194.420 14.670 195.970 14.890 ;
        RECT 196.350 14.880 196.780 14.940 ;
        RECT 197.160 14.890 197.610 14.940 ;
        RECT 198.210 14.890 198.710 15.280 ;
        RECT 197.160 14.670 198.710 14.890 ;
        RECT 207.920 15.280 209.470 15.500 ;
        RECT 207.920 14.890 208.420 15.280 ;
        RECT 209.020 15.230 209.470 15.280 ;
        RECT 209.850 15.230 210.280 15.290 ;
        RECT 210.660 15.280 212.210 15.500 ;
        RECT 214.960 15.430 215.370 15.860 ;
        RECT 215.760 15.760 216.210 15.860 ;
        RECT 210.660 15.230 211.110 15.280 ;
        RECT 209.020 14.940 211.110 15.230 ;
        RECT 209.020 14.890 209.470 14.940 ;
        RECT 192.270 14.310 192.720 14.380 ;
        RECT 190.420 14.070 192.720 14.310 ;
        RECT 190.420 13.960 190.870 14.070 ;
        RECT 192.270 13.960 192.720 14.070 ;
        RECT 193.670 14.310 194.120 14.410 ;
        RECT 195.520 14.310 195.970 14.410 ;
        RECT 193.670 14.070 195.970 14.310 ;
        RECT 193.670 13.990 194.120 14.070 ;
        RECT 174.180 13.410 175.710 13.620 ;
        RECT 176.090 13.410 176.540 13.500 ;
        RECT 176.920 13.410 178.450 13.620 ;
        RECT 187.680 13.620 188.130 13.900 ;
        RECT 191.500 13.620 191.950 13.900 ;
        RECT 194.720 13.630 195.130 14.070 ;
        RECT 195.520 13.960 195.970 14.070 ;
        RECT 197.160 14.310 197.610 14.410 ;
        RECT 199.010 14.310 199.460 14.410 ;
        RECT 197.160 14.070 199.460 14.310 ;
        RECT 197.160 13.960 197.610 14.070 ;
        RECT 198.000 13.630 198.410 14.070 ;
        RECT 199.010 13.990 199.460 14.070 ;
        RECT 200.410 14.310 200.860 14.380 ;
        RECT 201.460 14.310 201.870 14.740 ;
        RECT 202.260 14.310 202.710 14.410 ;
        RECT 200.410 14.070 202.710 14.310 ;
        RECT 200.410 13.960 200.860 14.070 ;
        RECT 202.260 13.960 202.710 14.070 ;
        RECT 203.920 14.310 204.370 14.410 ;
        RECT 204.760 14.310 205.170 14.740 ;
        RECT 207.920 14.670 209.470 14.890 ;
        RECT 209.850 14.880 210.280 14.940 ;
        RECT 210.660 14.890 211.110 14.940 ;
        RECT 211.710 14.890 212.210 15.280 ;
        RECT 210.660 14.670 212.210 14.890 ;
        RECT 205.770 14.310 206.220 14.380 ;
        RECT 203.920 14.070 206.220 14.310 ;
        RECT 203.920 13.960 204.370 14.070 ;
        RECT 205.770 13.960 206.220 14.070 ;
        RECT 207.170 14.310 207.620 14.410 ;
        RECT 209.020 14.310 209.470 14.410 ;
        RECT 207.170 14.070 209.470 14.310 ;
        RECT 207.170 13.990 207.620 14.070 ;
        RECT 187.680 13.410 189.210 13.620 ;
        RECT 189.590 13.410 190.040 13.500 ;
        RECT 190.420 13.410 191.950 13.620 ;
        RECT 201.180 13.620 201.630 13.900 ;
        RECT 205.000 13.620 205.450 13.900 ;
        RECT 208.220 13.630 208.630 14.070 ;
        RECT 209.020 13.960 209.470 14.070 ;
        RECT 210.660 14.310 211.110 14.410 ;
        RECT 212.510 14.310 212.960 14.410 ;
        RECT 210.660 14.070 212.960 14.310 ;
        RECT 210.660 13.960 211.110 14.070 ;
        RECT 211.500 13.630 211.910 14.070 ;
        RECT 212.510 13.990 212.960 14.070 ;
        RECT 213.910 14.310 214.360 14.380 ;
        RECT 214.960 14.310 215.370 14.740 ;
        RECT 215.760 14.310 216.210 14.410 ;
        RECT 213.910 14.070 216.210 14.310 ;
        RECT 213.910 13.960 214.360 14.070 ;
        RECT 215.760 13.960 216.210 14.070 ;
        RECT 201.180 13.410 202.710 13.620 ;
        RECT 203.090 13.410 203.540 13.500 ;
        RECT 203.920 13.410 205.450 13.620 ;
        RECT 214.680 13.620 215.130 13.900 ;
        RECT 214.680 13.410 216.210 13.620 ;
        RECT 216.590 13.410 217.030 13.500 ;
        RECT 13.260 13.150 15.370 13.410 ;
        RECT 26.760 13.150 28.870 13.410 ;
        RECT 40.260 13.150 42.370 13.410 ;
        RECT 53.760 13.150 55.870 13.410 ;
        RECT 67.260 13.150 69.370 13.410 ;
        RECT 80.760 13.150 82.870 13.410 ;
        RECT 94.260 13.150 96.370 13.410 ;
        RECT 107.760 13.150 109.870 13.410 ;
        RECT 121.260 13.150 123.370 13.410 ;
        RECT 134.760 13.150 136.870 13.410 ;
        RECT 148.260 13.150 150.370 13.410 ;
        RECT 161.760 13.150 163.870 13.410 ;
        RECT 175.260 13.150 177.370 13.410 ;
        RECT 188.760 13.150 190.870 13.410 ;
        RECT 202.260 13.150 204.370 13.410 ;
        RECT 215.760 13.400 217.030 13.410 ;
        RECT 215.760 13.210 217.240 13.400 ;
        RECT 215.760 13.150 217.030 13.210 ;
        RECT 12.180 12.940 13.710 13.150 ;
        RECT 14.090 13.060 14.540 13.150 ;
        RECT 14.920 12.940 16.450 13.150 ;
        RECT 1.420 12.490 1.870 12.600 ;
        RECT 3.270 12.490 3.720 12.600 ;
        RECT 1.420 12.250 3.720 12.490 ;
        RECT 1.420 12.150 1.870 12.250 ;
        RECT 2.260 11.820 2.670 12.250 ;
        RECT 3.270 12.180 3.720 12.250 ;
        RECT 4.670 12.490 5.120 12.570 ;
        RECT 5.720 12.490 6.130 12.930 ;
        RECT 6.520 12.490 6.970 12.600 ;
        RECT 4.670 12.250 6.970 12.490 ;
        RECT 4.670 12.150 5.120 12.250 ;
        RECT 6.520 12.150 6.970 12.250 ;
        RECT 8.160 12.490 8.610 12.600 ;
        RECT 9.000 12.490 9.410 12.930 ;
        RECT 12.180 12.660 12.630 12.940 ;
        RECT 16.000 12.660 16.450 12.940 ;
        RECT 25.680 12.940 27.210 13.150 ;
        RECT 27.590 13.060 28.040 13.150 ;
        RECT 28.420 12.940 29.950 13.150 ;
        RECT 10.010 12.490 10.460 12.570 ;
        RECT 8.160 12.250 10.460 12.490 ;
        RECT 8.160 12.150 8.610 12.250 ;
        RECT 10.010 12.150 10.460 12.250 ;
        RECT 11.410 12.490 11.860 12.600 ;
        RECT 13.260 12.490 13.710 12.600 ;
        RECT 11.410 12.250 13.710 12.490 ;
        RECT 11.410 12.180 11.860 12.250 ;
        RECT 5.420 11.670 6.970 11.890 ;
        RECT 5.420 11.280 5.920 11.670 ;
        RECT 6.520 11.620 6.970 11.670 ;
        RECT 7.350 11.620 7.780 11.680 ;
        RECT 8.160 11.670 9.710 11.890 ;
        RECT 12.460 11.820 12.870 12.250 ;
        RECT 13.260 12.150 13.710 12.250 ;
        RECT 14.920 12.490 15.370 12.600 ;
        RECT 16.770 12.490 17.220 12.600 ;
        RECT 14.920 12.250 17.220 12.490 ;
        RECT 14.920 12.150 15.370 12.250 ;
        RECT 15.760 11.820 16.170 12.250 ;
        RECT 16.770 12.180 17.220 12.250 ;
        RECT 18.170 12.490 18.620 12.570 ;
        RECT 19.220 12.490 19.630 12.930 ;
        RECT 20.020 12.490 20.470 12.600 ;
        RECT 18.170 12.250 20.470 12.490 ;
        RECT 18.170 12.150 18.620 12.250 ;
        RECT 20.020 12.150 20.470 12.250 ;
        RECT 21.660 12.490 22.110 12.600 ;
        RECT 22.500 12.490 22.910 12.930 ;
        RECT 25.680 12.660 26.130 12.940 ;
        RECT 29.500 12.660 29.950 12.940 ;
        RECT 39.180 12.940 40.710 13.150 ;
        RECT 41.090 13.060 41.540 13.150 ;
        RECT 41.920 12.940 43.450 13.150 ;
        RECT 23.510 12.490 23.960 12.570 ;
        RECT 21.660 12.250 23.960 12.490 ;
        RECT 21.660 12.150 22.110 12.250 ;
        RECT 23.510 12.150 23.960 12.250 ;
        RECT 24.910 12.490 25.360 12.600 ;
        RECT 26.760 12.490 27.210 12.600 ;
        RECT 24.910 12.250 27.210 12.490 ;
        RECT 24.910 12.180 25.360 12.250 ;
        RECT 8.160 11.620 8.610 11.670 ;
        RECT 6.520 11.330 8.610 11.620 ;
        RECT 6.520 11.280 6.970 11.330 ;
        RECT 1.420 10.700 1.870 10.800 ;
        RECT 2.260 10.700 2.670 11.130 ;
        RECT 5.420 11.060 6.970 11.280 ;
        RECT 7.350 11.270 7.780 11.330 ;
        RECT 8.160 11.280 8.610 11.330 ;
        RECT 9.210 11.280 9.710 11.670 ;
        RECT 8.160 11.060 9.710 11.280 ;
        RECT 18.920 11.670 20.470 11.890 ;
        RECT 18.920 11.280 19.420 11.670 ;
        RECT 20.020 11.620 20.470 11.670 ;
        RECT 20.850 11.620 21.280 11.680 ;
        RECT 21.660 11.670 23.210 11.890 ;
        RECT 25.960 11.820 26.370 12.250 ;
        RECT 26.760 12.150 27.210 12.250 ;
        RECT 28.420 12.490 28.870 12.600 ;
        RECT 30.270 12.490 30.720 12.600 ;
        RECT 28.420 12.250 30.720 12.490 ;
        RECT 28.420 12.150 28.870 12.250 ;
        RECT 29.260 11.820 29.670 12.250 ;
        RECT 30.270 12.180 30.720 12.250 ;
        RECT 31.670 12.490 32.120 12.570 ;
        RECT 32.720 12.490 33.130 12.930 ;
        RECT 33.520 12.490 33.970 12.600 ;
        RECT 31.670 12.250 33.970 12.490 ;
        RECT 31.670 12.150 32.120 12.250 ;
        RECT 33.520 12.150 33.970 12.250 ;
        RECT 35.160 12.490 35.610 12.600 ;
        RECT 36.000 12.490 36.410 12.930 ;
        RECT 39.180 12.660 39.630 12.940 ;
        RECT 43.000 12.660 43.450 12.940 ;
        RECT 52.680 12.940 54.210 13.150 ;
        RECT 54.590 13.060 55.040 13.150 ;
        RECT 55.420 12.940 56.950 13.150 ;
        RECT 37.010 12.490 37.460 12.570 ;
        RECT 35.160 12.250 37.460 12.490 ;
        RECT 35.160 12.150 35.610 12.250 ;
        RECT 37.010 12.150 37.460 12.250 ;
        RECT 38.410 12.490 38.860 12.600 ;
        RECT 40.260 12.490 40.710 12.600 ;
        RECT 38.410 12.250 40.710 12.490 ;
        RECT 38.410 12.180 38.860 12.250 ;
        RECT 21.660 11.620 22.110 11.670 ;
        RECT 20.020 11.330 22.110 11.620 ;
        RECT 20.020 11.280 20.470 11.330 ;
        RECT 3.270 10.700 3.720 10.770 ;
        RECT 1.420 10.460 3.720 10.700 ;
        RECT 1.420 10.350 1.870 10.460 ;
        RECT 3.270 10.350 3.720 10.460 ;
        RECT 4.670 10.700 5.120 10.800 ;
        RECT 6.520 10.700 6.970 10.800 ;
        RECT 4.670 10.460 6.970 10.700 ;
        RECT 4.670 10.380 5.120 10.460 ;
        RECT 5.720 10.020 6.130 10.460 ;
        RECT 6.520 10.350 6.970 10.460 ;
        RECT 8.160 10.700 8.610 10.800 ;
        RECT 10.010 10.700 10.460 10.800 ;
        RECT 8.160 10.460 10.460 10.700 ;
        RECT 8.160 10.350 8.610 10.460 ;
        RECT 9.000 10.020 9.410 10.460 ;
        RECT 10.010 10.380 10.460 10.460 ;
        RECT 11.410 10.700 11.860 10.770 ;
        RECT 12.460 10.700 12.870 11.130 ;
        RECT 13.260 10.700 13.710 10.800 ;
        RECT 11.410 10.460 13.710 10.700 ;
        RECT 11.410 10.350 11.860 10.460 ;
        RECT 13.260 10.350 13.710 10.460 ;
        RECT 14.920 10.700 15.370 10.800 ;
        RECT 15.760 10.700 16.170 11.130 ;
        RECT 18.920 11.060 20.470 11.280 ;
        RECT 20.850 11.270 21.280 11.330 ;
        RECT 21.660 11.280 22.110 11.330 ;
        RECT 22.710 11.280 23.210 11.670 ;
        RECT 21.660 11.060 23.210 11.280 ;
        RECT 32.420 11.670 33.970 11.890 ;
        RECT 32.420 11.280 32.920 11.670 ;
        RECT 33.520 11.620 33.970 11.670 ;
        RECT 34.350 11.620 34.780 11.680 ;
        RECT 35.160 11.670 36.710 11.890 ;
        RECT 39.460 11.820 39.870 12.250 ;
        RECT 40.260 12.150 40.710 12.250 ;
        RECT 41.920 12.490 42.370 12.600 ;
        RECT 43.770 12.490 44.220 12.600 ;
        RECT 41.920 12.250 44.220 12.490 ;
        RECT 41.920 12.150 42.370 12.250 ;
        RECT 42.760 11.820 43.170 12.250 ;
        RECT 43.770 12.180 44.220 12.250 ;
        RECT 45.170 12.490 45.620 12.570 ;
        RECT 46.220 12.490 46.630 12.930 ;
        RECT 47.020 12.490 47.470 12.600 ;
        RECT 45.170 12.250 47.470 12.490 ;
        RECT 45.170 12.150 45.620 12.250 ;
        RECT 47.020 12.150 47.470 12.250 ;
        RECT 48.660 12.490 49.110 12.600 ;
        RECT 49.500 12.490 49.910 12.930 ;
        RECT 52.680 12.660 53.130 12.940 ;
        RECT 56.500 12.660 56.950 12.940 ;
        RECT 66.180 12.940 67.710 13.150 ;
        RECT 68.090 13.060 68.540 13.150 ;
        RECT 68.920 12.940 70.450 13.150 ;
        RECT 50.510 12.490 50.960 12.570 ;
        RECT 48.660 12.250 50.960 12.490 ;
        RECT 48.660 12.150 49.110 12.250 ;
        RECT 50.510 12.150 50.960 12.250 ;
        RECT 51.910 12.490 52.360 12.600 ;
        RECT 53.760 12.490 54.210 12.600 ;
        RECT 51.910 12.250 54.210 12.490 ;
        RECT 51.910 12.180 52.360 12.250 ;
        RECT 35.160 11.620 35.610 11.670 ;
        RECT 33.520 11.330 35.610 11.620 ;
        RECT 33.520 11.280 33.970 11.330 ;
        RECT 16.770 10.700 17.220 10.770 ;
        RECT 14.920 10.460 17.220 10.700 ;
        RECT 14.920 10.350 15.370 10.460 ;
        RECT 16.770 10.350 17.220 10.460 ;
        RECT 18.170 10.700 18.620 10.800 ;
        RECT 20.020 10.700 20.470 10.800 ;
        RECT 18.170 10.460 20.470 10.700 ;
        RECT 18.170 10.380 18.620 10.460 ;
        RECT 12.180 10.010 12.630 10.290 ;
        RECT 16.000 10.010 16.450 10.290 ;
        RECT 19.220 10.020 19.630 10.460 ;
        RECT 20.020 10.350 20.470 10.460 ;
        RECT 21.660 10.700 22.110 10.800 ;
        RECT 23.510 10.700 23.960 10.800 ;
        RECT 21.660 10.460 23.960 10.700 ;
        RECT 21.660 10.350 22.110 10.460 ;
        RECT 22.500 10.020 22.910 10.460 ;
        RECT 23.510 10.380 23.960 10.460 ;
        RECT 24.910 10.700 25.360 10.770 ;
        RECT 25.960 10.700 26.370 11.130 ;
        RECT 26.760 10.700 27.210 10.800 ;
        RECT 24.910 10.460 27.210 10.700 ;
        RECT 24.910 10.350 25.360 10.460 ;
        RECT 26.760 10.350 27.210 10.460 ;
        RECT 28.420 10.700 28.870 10.800 ;
        RECT 29.260 10.700 29.670 11.130 ;
        RECT 32.420 11.060 33.970 11.280 ;
        RECT 34.350 11.270 34.780 11.330 ;
        RECT 35.160 11.280 35.610 11.330 ;
        RECT 36.210 11.280 36.710 11.670 ;
        RECT 35.160 11.060 36.710 11.280 ;
        RECT 45.920 11.670 47.470 11.890 ;
        RECT 45.920 11.280 46.420 11.670 ;
        RECT 47.020 11.620 47.470 11.670 ;
        RECT 47.850 11.620 48.280 11.680 ;
        RECT 48.660 11.670 50.210 11.890 ;
        RECT 52.960 11.820 53.370 12.250 ;
        RECT 53.760 12.150 54.210 12.250 ;
        RECT 55.420 12.490 55.870 12.600 ;
        RECT 57.270 12.490 57.720 12.600 ;
        RECT 55.420 12.250 57.720 12.490 ;
        RECT 55.420 12.150 55.870 12.250 ;
        RECT 56.260 11.820 56.670 12.250 ;
        RECT 57.270 12.180 57.720 12.250 ;
        RECT 58.670 12.490 59.120 12.570 ;
        RECT 59.720 12.490 60.130 12.930 ;
        RECT 60.520 12.490 60.970 12.600 ;
        RECT 58.670 12.250 60.970 12.490 ;
        RECT 58.670 12.150 59.120 12.250 ;
        RECT 60.520 12.150 60.970 12.250 ;
        RECT 62.160 12.490 62.610 12.600 ;
        RECT 63.000 12.490 63.410 12.930 ;
        RECT 66.180 12.660 66.630 12.940 ;
        RECT 70.000 12.660 70.450 12.940 ;
        RECT 79.680 12.940 81.210 13.150 ;
        RECT 81.590 13.060 82.040 13.150 ;
        RECT 82.420 12.940 83.950 13.150 ;
        RECT 64.010 12.490 64.460 12.570 ;
        RECT 62.160 12.250 64.460 12.490 ;
        RECT 62.160 12.150 62.610 12.250 ;
        RECT 64.010 12.150 64.460 12.250 ;
        RECT 65.410 12.490 65.860 12.600 ;
        RECT 67.260 12.490 67.710 12.600 ;
        RECT 65.410 12.250 67.710 12.490 ;
        RECT 65.410 12.180 65.860 12.250 ;
        RECT 48.660 11.620 49.110 11.670 ;
        RECT 47.020 11.330 49.110 11.620 ;
        RECT 47.020 11.280 47.470 11.330 ;
        RECT 30.270 10.700 30.720 10.770 ;
        RECT 28.420 10.460 30.720 10.700 ;
        RECT 28.420 10.350 28.870 10.460 ;
        RECT 30.270 10.350 30.720 10.460 ;
        RECT 31.670 10.700 32.120 10.800 ;
        RECT 33.520 10.700 33.970 10.800 ;
        RECT 31.670 10.460 33.970 10.700 ;
        RECT 31.670 10.380 32.120 10.460 ;
        RECT 12.180 9.800 13.710 10.010 ;
        RECT 14.090 9.800 14.540 9.890 ;
        RECT 14.920 9.800 16.450 10.010 ;
        RECT 25.680 10.010 26.130 10.290 ;
        RECT 29.500 10.010 29.950 10.290 ;
        RECT 32.720 10.020 33.130 10.460 ;
        RECT 33.520 10.350 33.970 10.460 ;
        RECT 35.160 10.700 35.610 10.800 ;
        RECT 37.010 10.700 37.460 10.800 ;
        RECT 35.160 10.460 37.460 10.700 ;
        RECT 35.160 10.350 35.610 10.460 ;
        RECT 36.000 10.020 36.410 10.460 ;
        RECT 37.010 10.380 37.460 10.460 ;
        RECT 38.410 10.700 38.860 10.770 ;
        RECT 39.460 10.700 39.870 11.130 ;
        RECT 40.260 10.700 40.710 10.800 ;
        RECT 38.410 10.460 40.710 10.700 ;
        RECT 38.410 10.350 38.860 10.460 ;
        RECT 40.260 10.350 40.710 10.460 ;
        RECT 41.920 10.700 42.370 10.800 ;
        RECT 42.760 10.700 43.170 11.130 ;
        RECT 45.920 11.060 47.470 11.280 ;
        RECT 47.850 11.270 48.280 11.330 ;
        RECT 48.660 11.280 49.110 11.330 ;
        RECT 49.710 11.280 50.210 11.670 ;
        RECT 48.660 11.060 50.210 11.280 ;
        RECT 59.420 11.670 60.970 11.890 ;
        RECT 59.420 11.280 59.920 11.670 ;
        RECT 60.520 11.620 60.970 11.670 ;
        RECT 61.350 11.620 61.780 11.680 ;
        RECT 62.160 11.670 63.710 11.890 ;
        RECT 66.460 11.820 66.870 12.250 ;
        RECT 67.260 12.150 67.710 12.250 ;
        RECT 68.920 12.490 69.370 12.600 ;
        RECT 70.770 12.490 71.220 12.600 ;
        RECT 68.920 12.250 71.220 12.490 ;
        RECT 68.920 12.150 69.370 12.250 ;
        RECT 69.760 11.820 70.170 12.250 ;
        RECT 70.770 12.180 71.220 12.250 ;
        RECT 72.170 12.490 72.620 12.570 ;
        RECT 73.220 12.490 73.630 12.930 ;
        RECT 74.020 12.490 74.470 12.600 ;
        RECT 72.170 12.250 74.470 12.490 ;
        RECT 72.170 12.150 72.620 12.250 ;
        RECT 74.020 12.150 74.470 12.250 ;
        RECT 75.660 12.490 76.110 12.600 ;
        RECT 76.500 12.490 76.910 12.930 ;
        RECT 79.680 12.660 80.130 12.940 ;
        RECT 83.500 12.660 83.950 12.940 ;
        RECT 93.180 12.940 94.710 13.150 ;
        RECT 95.090 13.060 95.540 13.150 ;
        RECT 95.920 12.940 97.450 13.150 ;
        RECT 77.510 12.490 77.960 12.570 ;
        RECT 75.660 12.250 77.960 12.490 ;
        RECT 75.660 12.150 76.110 12.250 ;
        RECT 77.510 12.150 77.960 12.250 ;
        RECT 78.910 12.490 79.360 12.600 ;
        RECT 80.760 12.490 81.210 12.600 ;
        RECT 78.910 12.250 81.210 12.490 ;
        RECT 78.910 12.180 79.360 12.250 ;
        RECT 62.160 11.620 62.610 11.670 ;
        RECT 60.520 11.330 62.610 11.620 ;
        RECT 60.520 11.280 60.970 11.330 ;
        RECT 43.770 10.700 44.220 10.770 ;
        RECT 41.920 10.460 44.220 10.700 ;
        RECT 41.920 10.350 42.370 10.460 ;
        RECT 43.770 10.350 44.220 10.460 ;
        RECT 45.170 10.700 45.620 10.800 ;
        RECT 47.020 10.700 47.470 10.800 ;
        RECT 45.170 10.460 47.470 10.700 ;
        RECT 45.170 10.380 45.620 10.460 ;
        RECT 25.680 9.800 27.210 10.010 ;
        RECT 27.590 9.800 28.040 9.890 ;
        RECT 28.420 9.800 29.950 10.010 ;
        RECT 39.180 10.010 39.630 10.290 ;
        RECT 43.000 10.010 43.450 10.290 ;
        RECT 46.220 10.020 46.630 10.460 ;
        RECT 47.020 10.350 47.470 10.460 ;
        RECT 48.660 10.700 49.110 10.800 ;
        RECT 50.510 10.700 50.960 10.800 ;
        RECT 48.660 10.460 50.960 10.700 ;
        RECT 48.660 10.350 49.110 10.460 ;
        RECT 49.500 10.020 49.910 10.460 ;
        RECT 50.510 10.380 50.960 10.460 ;
        RECT 51.910 10.700 52.360 10.770 ;
        RECT 52.960 10.700 53.370 11.130 ;
        RECT 53.760 10.700 54.210 10.800 ;
        RECT 51.910 10.460 54.210 10.700 ;
        RECT 51.910 10.350 52.360 10.460 ;
        RECT 53.760 10.350 54.210 10.460 ;
        RECT 55.420 10.700 55.870 10.800 ;
        RECT 56.260 10.700 56.670 11.130 ;
        RECT 59.420 11.060 60.970 11.280 ;
        RECT 61.350 11.270 61.780 11.330 ;
        RECT 62.160 11.280 62.610 11.330 ;
        RECT 63.210 11.280 63.710 11.670 ;
        RECT 62.160 11.060 63.710 11.280 ;
        RECT 72.920 11.670 74.470 11.890 ;
        RECT 72.920 11.280 73.420 11.670 ;
        RECT 74.020 11.620 74.470 11.670 ;
        RECT 74.850 11.620 75.280 11.680 ;
        RECT 75.660 11.670 77.210 11.890 ;
        RECT 79.960 11.820 80.370 12.250 ;
        RECT 80.760 12.150 81.210 12.250 ;
        RECT 82.420 12.490 82.870 12.600 ;
        RECT 84.270 12.490 84.720 12.600 ;
        RECT 82.420 12.250 84.720 12.490 ;
        RECT 82.420 12.150 82.870 12.250 ;
        RECT 83.260 11.820 83.670 12.250 ;
        RECT 84.270 12.180 84.720 12.250 ;
        RECT 85.670 12.490 86.120 12.570 ;
        RECT 86.720 12.490 87.130 12.930 ;
        RECT 87.520 12.490 87.970 12.600 ;
        RECT 85.670 12.250 87.970 12.490 ;
        RECT 85.670 12.150 86.120 12.250 ;
        RECT 87.520 12.150 87.970 12.250 ;
        RECT 89.160 12.490 89.610 12.600 ;
        RECT 90.000 12.490 90.410 12.930 ;
        RECT 93.180 12.660 93.630 12.940 ;
        RECT 97.000 12.660 97.450 12.940 ;
        RECT 106.680 12.940 108.210 13.150 ;
        RECT 108.590 13.060 109.040 13.150 ;
        RECT 109.420 12.940 110.950 13.150 ;
        RECT 91.010 12.490 91.460 12.570 ;
        RECT 89.160 12.250 91.460 12.490 ;
        RECT 89.160 12.150 89.610 12.250 ;
        RECT 91.010 12.150 91.460 12.250 ;
        RECT 92.410 12.490 92.860 12.600 ;
        RECT 94.260 12.490 94.710 12.600 ;
        RECT 92.410 12.250 94.710 12.490 ;
        RECT 92.410 12.180 92.860 12.250 ;
        RECT 75.660 11.620 76.110 11.670 ;
        RECT 74.020 11.330 76.110 11.620 ;
        RECT 74.020 11.280 74.470 11.330 ;
        RECT 57.270 10.700 57.720 10.770 ;
        RECT 55.420 10.460 57.720 10.700 ;
        RECT 55.420 10.350 55.870 10.460 ;
        RECT 57.270 10.350 57.720 10.460 ;
        RECT 58.670 10.700 59.120 10.800 ;
        RECT 60.520 10.700 60.970 10.800 ;
        RECT 58.670 10.460 60.970 10.700 ;
        RECT 58.670 10.380 59.120 10.460 ;
        RECT 39.180 9.800 40.710 10.010 ;
        RECT 41.090 9.800 41.540 9.890 ;
        RECT 41.920 9.800 43.450 10.010 ;
        RECT 52.680 10.010 53.130 10.290 ;
        RECT 56.500 10.010 56.950 10.290 ;
        RECT 59.720 10.020 60.130 10.460 ;
        RECT 60.520 10.350 60.970 10.460 ;
        RECT 62.160 10.700 62.610 10.800 ;
        RECT 64.010 10.700 64.460 10.800 ;
        RECT 62.160 10.460 64.460 10.700 ;
        RECT 62.160 10.350 62.610 10.460 ;
        RECT 63.000 10.020 63.410 10.460 ;
        RECT 64.010 10.380 64.460 10.460 ;
        RECT 65.410 10.700 65.860 10.770 ;
        RECT 66.460 10.700 66.870 11.130 ;
        RECT 67.260 10.700 67.710 10.800 ;
        RECT 65.410 10.460 67.710 10.700 ;
        RECT 65.410 10.350 65.860 10.460 ;
        RECT 67.260 10.350 67.710 10.460 ;
        RECT 68.920 10.700 69.370 10.800 ;
        RECT 69.760 10.700 70.170 11.130 ;
        RECT 72.920 11.060 74.470 11.280 ;
        RECT 74.850 11.270 75.280 11.330 ;
        RECT 75.660 11.280 76.110 11.330 ;
        RECT 76.710 11.280 77.210 11.670 ;
        RECT 75.660 11.060 77.210 11.280 ;
        RECT 86.420 11.670 87.970 11.890 ;
        RECT 86.420 11.280 86.920 11.670 ;
        RECT 87.520 11.620 87.970 11.670 ;
        RECT 88.350 11.620 88.780 11.680 ;
        RECT 89.160 11.670 90.710 11.890 ;
        RECT 93.460 11.820 93.870 12.250 ;
        RECT 94.260 12.150 94.710 12.250 ;
        RECT 95.920 12.490 96.370 12.600 ;
        RECT 97.770 12.490 98.220 12.600 ;
        RECT 95.920 12.250 98.220 12.490 ;
        RECT 95.920 12.150 96.370 12.250 ;
        RECT 96.760 11.820 97.170 12.250 ;
        RECT 97.770 12.180 98.220 12.250 ;
        RECT 99.170 12.490 99.620 12.570 ;
        RECT 100.220 12.490 100.630 12.930 ;
        RECT 101.020 12.490 101.470 12.600 ;
        RECT 99.170 12.250 101.470 12.490 ;
        RECT 99.170 12.150 99.620 12.250 ;
        RECT 101.020 12.150 101.470 12.250 ;
        RECT 102.660 12.490 103.110 12.600 ;
        RECT 103.500 12.490 103.910 12.930 ;
        RECT 106.680 12.660 107.130 12.940 ;
        RECT 110.500 12.660 110.950 12.940 ;
        RECT 120.180 12.940 121.710 13.150 ;
        RECT 122.090 13.060 122.540 13.150 ;
        RECT 122.920 12.940 124.450 13.150 ;
        RECT 104.510 12.490 104.960 12.570 ;
        RECT 102.660 12.250 104.960 12.490 ;
        RECT 102.660 12.150 103.110 12.250 ;
        RECT 104.510 12.150 104.960 12.250 ;
        RECT 105.910 12.490 106.360 12.600 ;
        RECT 107.760 12.490 108.210 12.600 ;
        RECT 105.910 12.250 108.210 12.490 ;
        RECT 105.910 12.180 106.360 12.250 ;
        RECT 89.160 11.620 89.610 11.670 ;
        RECT 87.520 11.330 89.610 11.620 ;
        RECT 87.520 11.280 87.970 11.330 ;
        RECT 70.770 10.700 71.220 10.770 ;
        RECT 68.920 10.460 71.220 10.700 ;
        RECT 68.920 10.350 69.370 10.460 ;
        RECT 70.770 10.350 71.220 10.460 ;
        RECT 72.170 10.700 72.620 10.800 ;
        RECT 74.020 10.700 74.470 10.800 ;
        RECT 72.170 10.460 74.470 10.700 ;
        RECT 72.170 10.380 72.620 10.460 ;
        RECT 52.680 9.800 54.210 10.010 ;
        RECT 54.590 9.800 55.040 9.890 ;
        RECT 55.420 9.800 56.950 10.010 ;
        RECT 66.180 10.010 66.630 10.290 ;
        RECT 70.000 10.010 70.450 10.290 ;
        RECT 73.220 10.020 73.630 10.460 ;
        RECT 74.020 10.350 74.470 10.460 ;
        RECT 75.660 10.700 76.110 10.800 ;
        RECT 77.510 10.700 77.960 10.800 ;
        RECT 75.660 10.460 77.960 10.700 ;
        RECT 75.660 10.350 76.110 10.460 ;
        RECT 76.500 10.020 76.910 10.460 ;
        RECT 77.510 10.380 77.960 10.460 ;
        RECT 78.910 10.700 79.360 10.770 ;
        RECT 79.960 10.700 80.370 11.130 ;
        RECT 80.760 10.700 81.210 10.800 ;
        RECT 78.910 10.460 81.210 10.700 ;
        RECT 78.910 10.350 79.360 10.460 ;
        RECT 80.760 10.350 81.210 10.460 ;
        RECT 82.420 10.700 82.870 10.800 ;
        RECT 83.260 10.700 83.670 11.130 ;
        RECT 86.420 11.060 87.970 11.280 ;
        RECT 88.350 11.270 88.780 11.330 ;
        RECT 89.160 11.280 89.610 11.330 ;
        RECT 90.210 11.280 90.710 11.670 ;
        RECT 89.160 11.060 90.710 11.280 ;
        RECT 99.920 11.670 101.470 11.890 ;
        RECT 99.920 11.280 100.420 11.670 ;
        RECT 101.020 11.620 101.470 11.670 ;
        RECT 101.850 11.620 102.280 11.680 ;
        RECT 102.660 11.670 104.210 11.890 ;
        RECT 106.960 11.820 107.370 12.250 ;
        RECT 107.760 12.150 108.210 12.250 ;
        RECT 109.420 12.490 109.870 12.600 ;
        RECT 111.270 12.490 111.720 12.600 ;
        RECT 109.420 12.250 111.720 12.490 ;
        RECT 109.420 12.150 109.870 12.250 ;
        RECT 110.260 11.820 110.670 12.250 ;
        RECT 111.270 12.180 111.720 12.250 ;
        RECT 112.670 12.490 113.120 12.570 ;
        RECT 113.720 12.490 114.130 12.930 ;
        RECT 114.520 12.490 114.970 12.600 ;
        RECT 112.670 12.250 114.970 12.490 ;
        RECT 112.670 12.150 113.120 12.250 ;
        RECT 114.520 12.150 114.970 12.250 ;
        RECT 116.160 12.490 116.610 12.600 ;
        RECT 117.000 12.490 117.410 12.930 ;
        RECT 120.180 12.660 120.630 12.940 ;
        RECT 124.000 12.660 124.450 12.940 ;
        RECT 133.680 12.940 135.210 13.150 ;
        RECT 135.590 13.060 136.040 13.150 ;
        RECT 136.420 12.940 137.950 13.150 ;
        RECT 118.010 12.490 118.460 12.570 ;
        RECT 116.160 12.250 118.460 12.490 ;
        RECT 116.160 12.150 116.610 12.250 ;
        RECT 118.010 12.150 118.460 12.250 ;
        RECT 119.410 12.490 119.860 12.600 ;
        RECT 121.260 12.490 121.710 12.600 ;
        RECT 119.410 12.250 121.710 12.490 ;
        RECT 119.410 12.180 119.860 12.250 ;
        RECT 102.660 11.620 103.110 11.670 ;
        RECT 101.020 11.330 103.110 11.620 ;
        RECT 101.020 11.280 101.470 11.330 ;
        RECT 84.270 10.700 84.720 10.770 ;
        RECT 82.420 10.460 84.720 10.700 ;
        RECT 82.420 10.350 82.870 10.460 ;
        RECT 84.270 10.350 84.720 10.460 ;
        RECT 85.670 10.700 86.120 10.800 ;
        RECT 87.520 10.700 87.970 10.800 ;
        RECT 85.670 10.460 87.970 10.700 ;
        RECT 85.670 10.380 86.120 10.460 ;
        RECT 66.180 9.800 67.710 10.010 ;
        RECT 68.090 9.800 68.540 9.890 ;
        RECT 68.920 9.800 70.450 10.010 ;
        RECT 79.680 10.010 80.130 10.290 ;
        RECT 83.500 10.010 83.950 10.290 ;
        RECT 86.720 10.020 87.130 10.460 ;
        RECT 87.520 10.350 87.970 10.460 ;
        RECT 89.160 10.700 89.610 10.800 ;
        RECT 91.010 10.700 91.460 10.800 ;
        RECT 89.160 10.460 91.460 10.700 ;
        RECT 89.160 10.350 89.610 10.460 ;
        RECT 90.000 10.020 90.410 10.460 ;
        RECT 91.010 10.380 91.460 10.460 ;
        RECT 92.410 10.700 92.860 10.770 ;
        RECT 93.460 10.700 93.870 11.130 ;
        RECT 94.260 10.700 94.710 10.800 ;
        RECT 92.410 10.460 94.710 10.700 ;
        RECT 92.410 10.350 92.860 10.460 ;
        RECT 94.260 10.350 94.710 10.460 ;
        RECT 95.920 10.700 96.370 10.800 ;
        RECT 96.760 10.700 97.170 11.130 ;
        RECT 99.920 11.060 101.470 11.280 ;
        RECT 101.850 11.270 102.280 11.330 ;
        RECT 102.660 11.280 103.110 11.330 ;
        RECT 103.710 11.280 104.210 11.670 ;
        RECT 102.660 11.060 104.210 11.280 ;
        RECT 113.420 11.670 114.970 11.890 ;
        RECT 113.420 11.280 113.920 11.670 ;
        RECT 114.520 11.620 114.970 11.670 ;
        RECT 115.350 11.620 115.780 11.680 ;
        RECT 116.160 11.670 117.710 11.890 ;
        RECT 120.460 11.820 120.870 12.250 ;
        RECT 121.260 12.150 121.710 12.250 ;
        RECT 122.920 12.490 123.370 12.600 ;
        RECT 124.770 12.490 125.220 12.600 ;
        RECT 122.920 12.250 125.220 12.490 ;
        RECT 122.920 12.150 123.370 12.250 ;
        RECT 123.760 11.820 124.170 12.250 ;
        RECT 124.770 12.180 125.220 12.250 ;
        RECT 126.170 12.490 126.620 12.570 ;
        RECT 127.220 12.490 127.630 12.930 ;
        RECT 128.020 12.490 128.470 12.600 ;
        RECT 126.170 12.250 128.470 12.490 ;
        RECT 126.170 12.150 126.620 12.250 ;
        RECT 128.020 12.150 128.470 12.250 ;
        RECT 129.660 12.490 130.110 12.600 ;
        RECT 130.500 12.490 130.910 12.930 ;
        RECT 133.680 12.660 134.130 12.940 ;
        RECT 137.500 12.660 137.950 12.940 ;
        RECT 147.180 12.940 148.710 13.150 ;
        RECT 149.090 13.060 149.540 13.150 ;
        RECT 149.920 12.940 151.450 13.150 ;
        RECT 131.510 12.490 131.960 12.570 ;
        RECT 129.660 12.250 131.960 12.490 ;
        RECT 129.660 12.150 130.110 12.250 ;
        RECT 131.510 12.150 131.960 12.250 ;
        RECT 132.910 12.490 133.360 12.600 ;
        RECT 134.760 12.490 135.210 12.600 ;
        RECT 132.910 12.250 135.210 12.490 ;
        RECT 132.910 12.180 133.360 12.250 ;
        RECT 116.160 11.620 116.610 11.670 ;
        RECT 114.520 11.330 116.610 11.620 ;
        RECT 114.520 11.280 114.970 11.330 ;
        RECT 97.770 10.700 98.220 10.770 ;
        RECT 95.920 10.460 98.220 10.700 ;
        RECT 95.920 10.350 96.370 10.460 ;
        RECT 97.770 10.350 98.220 10.460 ;
        RECT 99.170 10.700 99.620 10.800 ;
        RECT 101.020 10.700 101.470 10.800 ;
        RECT 99.170 10.460 101.470 10.700 ;
        RECT 99.170 10.380 99.620 10.460 ;
        RECT 79.680 9.800 81.210 10.010 ;
        RECT 81.590 9.800 82.040 9.890 ;
        RECT 82.420 9.800 83.950 10.010 ;
        RECT 93.180 10.010 93.630 10.290 ;
        RECT 97.000 10.010 97.450 10.290 ;
        RECT 100.220 10.020 100.630 10.460 ;
        RECT 101.020 10.350 101.470 10.460 ;
        RECT 102.660 10.700 103.110 10.800 ;
        RECT 104.510 10.700 104.960 10.800 ;
        RECT 102.660 10.460 104.960 10.700 ;
        RECT 102.660 10.350 103.110 10.460 ;
        RECT 103.500 10.020 103.910 10.460 ;
        RECT 104.510 10.380 104.960 10.460 ;
        RECT 105.910 10.700 106.360 10.770 ;
        RECT 106.960 10.700 107.370 11.130 ;
        RECT 107.760 10.700 108.210 10.800 ;
        RECT 105.910 10.460 108.210 10.700 ;
        RECT 105.910 10.350 106.360 10.460 ;
        RECT 107.760 10.350 108.210 10.460 ;
        RECT 109.420 10.700 109.870 10.800 ;
        RECT 110.260 10.700 110.670 11.130 ;
        RECT 113.420 11.060 114.970 11.280 ;
        RECT 115.350 11.270 115.780 11.330 ;
        RECT 116.160 11.280 116.610 11.330 ;
        RECT 117.210 11.280 117.710 11.670 ;
        RECT 116.160 11.060 117.710 11.280 ;
        RECT 126.920 11.670 128.470 11.890 ;
        RECT 126.920 11.280 127.420 11.670 ;
        RECT 128.020 11.620 128.470 11.670 ;
        RECT 128.850 11.620 129.280 11.680 ;
        RECT 129.660 11.670 131.210 11.890 ;
        RECT 133.960 11.820 134.370 12.250 ;
        RECT 134.760 12.150 135.210 12.250 ;
        RECT 136.420 12.490 136.870 12.600 ;
        RECT 138.270 12.490 138.720 12.600 ;
        RECT 136.420 12.250 138.720 12.490 ;
        RECT 136.420 12.150 136.870 12.250 ;
        RECT 137.260 11.820 137.670 12.250 ;
        RECT 138.270 12.180 138.720 12.250 ;
        RECT 139.670 12.490 140.120 12.570 ;
        RECT 140.720 12.490 141.130 12.930 ;
        RECT 141.520 12.490 141.970 12.600 ;
        RECT 139.670 12.250 141.970 12.490 ;
        RECT 139.670 12.150 140.120 12.250 ;
        RECT 141.520 12.150 141.970 12.250 ;
        RECT 143.160 12.490 143.610 12.600 ;
        RECT 144.000 12.490 144.410 12.930 ;
        RECT 147.180 12.660 147.630 12.940 ;
        RECT 151.000 12.660 151.450 12.940 ;
        RECT 160.680 12.940 162.210 13.150 ;
        RECT 162.590 13.060 163.040 13.150 ;
        RECT 163.420 12.940 164.950 13.150 ;
        RECT 145.010 12.490 145.460 12.570 ;
        RECT 143.160 12.250 145.460 12.490 ;
        RECT 143.160 12.150 143.610 12.250 ;
        RECT 145.010 12.150 145.460 12.250 ;
        RECT 146.410 12.490 146.860 12.600 ;
        RECT 148.260 12.490 148.710 12.600 ;
        RECT 146.410 12.250 148.710 12.490 ;
        RECT 146.410 12.180 146.860 12.250 ;
        RECT 129.660 11.620 130.110 11.670 ;
        RECT 128.020 11.330 130.110 11.620 ;
        RECT 128.020 11.280 128.470 11.330 ;
        RECT 111.270 10.700 111.720 10.770 ;
        RECT 109.420 10.460 111.720 10.700 ;
        RECT 109.420 10.350 109.870 10.460 ;
        RECT 111.270 10.350 111.720 10.460 ;
        RECT 112.670 10.700 113.120 10.800 ;
        RECT 114.520 10.700 114.970 10.800 ;
        RECT 112.670 10.460 114.970 10.700 ;
        RECT 112.670 10.380 113.120 10.460 ;
        RECT 93.180 9.800 94.710 10.010 ;
        RECT 95.090 9.800 95.540 9.890 ;
        RECT 95.920 9.800 97.450 10.010 ;
        RECT 106.680 10.010 107.130 10.290 ;
        RECT 110.500 10.010 110.950 10.290 ;
        RECT 113.720 10.020 114.130 10.460 ;
        RECT 114.520 10.350 114.970 10.460 ;
        RECT 116.160 10.700 116.610 10.800 ;
        RECT 118.010 10.700 118.460 10.800 ;
        RECT 116.160 10.460 118.460 10.700 ;
        RECT 116.160 10.350 116.610 10.460 ;
        RECT 117.000 10.020 117.410 10.460 ;
        RECT 118.010 10.380 118.460 10.460 ;
        RECT 119.410 10.700 119.860 10.770 ;
        RECT 120.460 10.700 120.870 11.130 ;
        RECT 121.260 10.700 121.710 10.800 ;
        RECT 119.410 10.460 121.710 10.700 ;
        RECT 119.410 10.350 119.860 10.460 ;
        RECT 121.260 10.350 121.710 10.460 ;
        RECT 122.920 10.700 123.370 10.800 ;
        RECT 123.760 10.700 124.170 11.130 ;
        RECT 126.920 11.060 128.470 11.280 ;
        RECT 128.850 11.270 129.280 11.330 ;
        RECT 129.660 11.280 130.110 11.330 ;
        RECT 130.710 11.280 131.210 11.670 ;
        RECT 129.660 11.060 131.210 11.280 ;
        RECT 140.420 11.670 141.970 11.890 ;
        RECT 140.420 11.280 140.920 11.670 ;
        RECT 141.520 11.620 141.970 11.670 ;
        RECT 142.350 11.620 142.780 11.680 ;
        RECT 143.160 11.670 144.710 11.890 ;
        RECT 147.460 11.820 147.870 12.250 ;
        RECT 148.260 12.150 148.710 12.250 ;
        RECT 149.920 12.490 150.370 12.600 ;
        RECT 151.770 12.490 152.220 12.600 ;
        RECT 149.920 12.250 152.220 12.490 ;
        RECT 149.920 12.150 150.370 12.250 ;
        RECT 150.760 11.820 151.170 12.250 ;
        RECT 151.770 12.180 152.220 12.250 ;
        RECT 153.170 12.490 153.620 12.570 ;
        RECT 154.220 12.490 154.630 12.930 ;
        RECT 155.020 12.490 155.470 12.600 ;
        RECT 153.170 12.250 155.470 12.490 ;
        RECT 153.170 12.150 153.620 12.250 ;
        RECT 155.020 12.150 155.470 12.250 ;
        RECT 156.660 12.490 157.110 12.600 ;
        RECT 157.500 12.490 157.910 12.930 ;
        RECT 160.680 12.660 161.130 12.940 ;
        RECT 164.500 12.660 164.950 12.940 ;
        RECT 174.180 12.940 175.710 13.150 ;
        RECT 176.090 13.060 176.540 13.150 ;
        RECT 176.920 12.940 178.450 13.150 ;
        RECT 158.510 12.490 158.960 12.570 ;
        RECT 156.660 12.250 158.960 12.490 ;
        RECT 156.660 12.150 157.110 12.250 ;
        RECT 158.510 12.150 158.960 12.250 ;
        RECT 159.910 12.490 160.360 12.600 ;
        RECT 161.760 12.490 162.210 12.600 ;
        RECT 159.910 12.250 162.210 12.490 ;
        RECT 159.910 12.180 160.360 12.250 ;
        RECT 143.160 11.620 143.610 11.670 ;
        RECT 141.520 11.330 143.610 11.620 ;
        RECT 141.520 11.280 141.970 11.330 ;
        RECT 124.770 10.700 125.220 10.770 ;
        RECT 122.920 10.460 125.220 10.700 ;
        RECT 122.920 10.350 123.370 10.460 ;
        RECT 124.770 10.350 125.220 10.460 ;
        RECT 126.170 10.700 126.620 10.800 ;
        RECT 128.020 10.700 128.470 10.800 ;
        RECT 126.170 10.460 128.470 10.700 ;
        RECT 126.170 10.380 126.620 10.460 ;
        RECT 106.680 9.800 108.210 10.010 ;
        RECT 108.590 9.800 109.040 9.890 ;
        RECT 109.420 9.800 110.950 10.010 ;
        RECT 120.180 10.010 120.630 10.290 ;
        RECT 124.000 10.010 124.450 10.290 ;
        RECT 127.220 10.020 127.630 10.460 ;
        RECT 128.020 10.350 128.470 10.460 ;
        RECT 129.660 10.700 130.110 10.800 ;
        RECT 131.510 10.700 131.960 10.800 ;
        RECT 129.660 10.460 131.960 10.700 ;
        RECT 129.660 10.350 130.110 10.460 ;
        RECT 130.500 10.020 130.910 10.460 ;
        RECT 131.510 10.380 131.960 10.460 ;
        RECT 132.910 10.700 133.360 10.770 ;
        RECT 133.960 10.700 134.370 11.130 ;
        RECT 134.760 10.700 135.210 10.800 ;
        RECT 132.910 10.460 135.210 10.700 ;
        RECT 132.910 10.350 133.360 10.460 ;
        RECT 134.760 10.350 135.210 10.460 ;
        RECT 136.420 10.700 136.870 10.800 ;
        RECT 137.260 10.700 137.670 11.130 ;
        RECT 140.420 11.060 141.970 11.280 ;
        RECT 142.350 11.270 142.780 11.330 ;
        RECT 143.160 11.280 143.610 11.330 ;
        RECT 144.210 11.280 144.710 11.670 ;
        RECT 143.160 11.060 144.710 11.280 ;
        RECT 153.920 11.670 155.470 11.890 ;
        RECT 153.920 11.280 154.420 11.670 ;
        RECT 155.020 11.620 155.470 11.670 ;
        RECT 155.850 11.620 156.280 11.680 ;
        RECT 156.660 11.670 158.210 11.890 ;
        RECT 160.960 11.820 161.370 12.250 ;
        RECT 161.760 12.150 162.210 12.250 ;
        RECT 163.420 12.490 163.870 12.600 ;
        RECT 165.270 12.490 165.720 12.600 ;
        RECT 163.420 12.250 165.720 12.490 ;
        RECT 163.420 12.150 163.870 12.250 ;
        RECT 164.260 11.820 164.670 12.250 ;
        RECT 165.270 12.180 165.720 12.250 ;
        RECT 166.670 12.490 167.120 12.570 ;
        RECT 167.720 12.490 168.130 12.930 ;
        RECT 168.520 12.490 168.970 12.600 ;
        RECT 166.670 12.250 168.970 12.490 ;
        RECT 166.670 12.150 167.120 12.250 ;
        RECT 168.520 12.150 168.970 12.250 ;
        RECT 170.160 12.490 170.610 12.600 ;
        RECT 171.000 12.490 171.410 12.930 ;
        RECT 174.180 12.660 174.630 12.940 ;
        RECT 178.000 12.660 178.450 12.940 ;
        RECT 187.680 12.940 189.210 13.150 ;
        RECT 189.590 13.060 190.040 13.150 ;
        RECT 190.420 12.940 191.950 13.150 ;
        RECT 172.010 12.490 172.460 12.570 ;
        RECT 170.160 12.250 172.460 12.490 ;
        RECT 170.160 12.150 170.610 12.250 ;
        RECT 172.010 12.150 172.460 12.250 ;
        RECT 173.410 12.490 173.860 12.600 ;
        RECT 175.260 12.490 175.710 12.600 ;
        RECT 173.410 12.250 175.710 12.490 ;
        RECT 173.410 12.180 173.860 12.250 ;
        RECT 156.660 11.620 157.110 11.670 ;
        RECT 155.020 11.330 157.110 11.620 ;
        RECT 155.020 11.280 155.470 11.330 ;
        RECT 138.270 10.700 138.720 10.770 ;
        RECT 136.420 10.460 138.720 10.700 ;
        RECT 136.420 10.350 136.870 10.460 ;
        RECT 138.270 10.350 138.720 10.460 ;
        RECT 139.670 10.700 140.120 10.800 ;
        RECT 141.520 10.700 141.970 10.800 ;
        RECT 139.670 10.460 141.970 10.700 ;
        RECT 139.670 10.380 140.120 10.460 ;
        RECT 120.180 9.800 121.710 10.010 ;
        RECT 122.090 9.800 122.540 9.890 ;
        RECT 122.920 9.800 124.450 10.010 ;
        RECT 133.680 10.010 134.130 10.290 ;
        RECT 137.500 10.010 137.950 10.290 ;
        RECT 140.720 10.020 141.130 10.460 ;
        RECT 141.520 10.350 141.970 10.460 ;
        RECT 143.160 10.700 143.610 10.800 ;
        RECT 145.010 10.700 145.460 10.800 ;
        RECT 143.160 10.460 145.460 10.700 ;
        RECT 143.160 10.350 143.610 10.460 ;
        RECT 144.000 10.020 144.410 10.460 ;
        RECT 145.010 10.380 145.460 10.460 ;
        RECT 146.410 10.700 146.860 10.770 ;
        RECT 147.460 10.700 147.870 11.130 ;
        RECT 148.260 10.700 148.710 10.800 ;
        RECT 146.410 10.460 148.710 10.700 ;
        RECT 146.410 10.350 146.860 10.460 ;
        RECT 148.260 10.350 148.710 10.460 ;
        RECT 149.920 10.700 150.370 10.800 ;
        RECT 150.760 10.700 151.170 11.130 ;
        RECT 153.920 11.060 155.470 11.280 ;
        RECT 155.850 11.270 156.280 11.330 ;
        RECT 156.660 11.280 157.110 11.330 ;
        RECT 157.710 11.280 158.210 11.670 ;
        RECT 156.660 11.060 158.210 11.280 ;
        RECT 167.420 11.670 168.970 11.890 ;
        RECT 167.420 11.280 167.920 11.670 ;
        RECT 168.520 11.620 168.970 11.670 ;
        RECT 169.350 11.620 169.780 11.680 ;
        RECT 170.160 11.670 171.710 11.890 ;
        RECT 174.460 11.820 174.870 12.250 ;
        RECT 175.260 12.150 175.710 12.250 ;
        RECT 176.920 12.490 177.370 12.600 ;
        RECT 178.770 12.490 179.220 12.600 ;
        RECT 176.920 12.250 179.220 12.490 ;
        RECT 176.920 12.150 177.370 12.250 ;
        RECT 177.760 11.820 178.170 12.250 ;
        RECT 178.770 12.180 179.220 12.250 ;
        RECT 180.170 12.490 180.620 12.570 ;
        RECT 181.220 12.490 181.630 12.930 ;
        RECT 182.020 12.490 182.470 12.600 ;
        RECT 180.170 12.250 182.470 12.490 ;
        RECT 180.170 12.150 180.620 12.250 ;
        RECT 182.020 12.150 182.470 12.250 ;
        RECT 183.660 12.490 184.110 12.600 ;
        RECT 184.500 12.490 184.910 12.930 ;
        RECT 187.680 12.660 188.130 12.940 ;
        RECT 191.500 12.660 191.950 12.940 ;
        RECT 201.180 12.940 202.710 13.150 ;
        RECT 203.090 13.060 203.540 13.150 ;
        RECT 203.920 12.940 205.450 13.150 ;
        RECT 185.510 12.490 185.960 12.570 ;
        RECT 183.660 12.250 185.960 12.490 ;
        RECT 183.660 12.150 184.110 12.250 ;
        RECT 185.510 12.150 185.960 12.250 ;
        RECT 186.910 12.490 187.360 12.600 ;
        RECT 188.760 12.490 189.210 12.600 ;
        RECT 186.910 12.250 189.210 12.490 ;
        RECT 186.910 12.180 187.360 12.250 ;
        RECT 170.160 11.620 170.610 11.670 ;
        RECT 168.520 11.330 170.610 11.620 ;
        RECT 168.520 11.280 168.970 11.330 ;
        RECT 151.770 10.700 152.220 10.770 ;
        RECT 149.920 10.460 152.220 10.700 ;
        RECT 149.920 10.350 150.370 10.460 ;
        RECT 151.770 10.350 152.220 10.460 ;
        RECT 153.170 10.700 153.620 10.800 ;
        RECT 155.020 10.700 155.470 10.800 ;
        RECT 153.170 10.460 155.470 10.700 ;
        RECT 153.170 10.380 153.620 10.460 ;
        RECT 133.680 9.800 135.210 10.010 ;
        RECT 135.590 9.800 136.040 9.890 ;
        RECT 136.420 9.800 137.950 10.010 ;
        RECT 147.180 10.010 147.630 10.290 ;
        RECT 151.000 10.010 151.450 10.290 ;
        RECT 154.220 10.020 154.630 10.460 ;
        RECT 155.020 10.350 155.470 10.460 ;
        RECT 156.660 10.700 157.110 10.800 ;
        RECT 158.510 10.700 158.960 10.800 ;
        RECT 156.660 10.460 158.960 10.700 ;
        RECT 156.660 10.350 157.110 10.460 ;
        RECT 157.500 10.020 157.910 10.460 ;
        RECT 158.510 10.380 158.960 10.460 ;
        RECT 159.910 10.700 160.360 10.770 ;
        RECT 160.960 10.700 161.370 11.130 ;
        RECT 161.760 10.700 162.210 10.800 ;
        RECT 159.910 10.460 162.210 10.700 ;
        RECT 159.910 10.350 160.360 10.460 ;
        RECT 161.760 10.350 162.210 10.460 ;
        RECT 163.420 10.700 163.870 10.800 ;
        RECT 164.260 10.700 164.670 11.130 ;
        RECT 167.420 11.060 168.970 11.280 ;
        RECT 169.350 11.270 169.780 11.330 ;
        RECT 170.160 11.280 170.610 11.330 ;
        RECT 171.210 11.280 171.710 11.670 ;
        RECT 170.160 11.060 171.710 11.280 ;
        RECT 180.920 11.670 182.470 11.890 ;
        RECT 180.920 11.280 181.420 11.670 ;
        RECT 182.020 11.620 182.470 11.670 ;
        RECT 182.850 11.620 183.280 11.680 ;
        RECT 183.660 11.670 185.210 11.890 ;
        RECT 187.960 11.820 188.370 12.250 ;
        RECT 188.760 12.150 189.210 12.250 ;
        RECT 190.420 12.490 190.870 12.600 ;
        RECT 192.270 12.490 192.720 12.600 ;
        RECT 190.420 12.250 192.720 12.490 ;
        RECT 190.420 12.150 190.870 12.250 ;
        RECT 191.260 11.820 191.670 12.250 ;
        RECT 192.270 12.180 192.720 12.250 ;
        RECT 193.670 12.490 194.120 12.570 ;
        RECT 194.720 12.490 195.130 12.930 ;
        RECT 195.520 12.490 195.970 12.600 ;
        RECT 193.670 12.250 195.970 12.490 ;
        RECT 193.670 12.150 194.120 12.250 ;
        RECT 195.520 12.150 195.970 12.250 ;
        RECT 197.160 12.490 197.610 12.600 ;
        RECT 198.000 12.490 198.410 12.930 ;
        RECT 201.180 12.660 201.630 12.940 ;
        RECT 205.000 12.660 205.450 12.940 ;
        RECT 214.680 12.940 216.210 13.150 ;
        RECT 216.590 13.060 217.030 13.150 ;
        RECT 199.010 12.490 199.460 12.570 ;
        RECT 197.160 12.250 199.460 12.490 ;
        RECT 197.160 12.150 197.610 12.250 ;
        RECT 199.010 12.150 199.460 12.250 ;
        RECT 200.410 12.490 200.860 12.600 ;
        RECT 202.260 12.490 202.710 12.600 ;
        RECT 200.410 12.250 202.710 12.490 ;
        RECT 200.410 12.180 200.860 12.250 ;
        RECT 183.660 11.620 184.110 11.670 ;
        RECT 182.020 11.330 184.110 11.620 ;
        RECT 182.020 11.280 182.470 11.330 ;
        RECT 165.270 10.700 165.720 10.770 ;
        RECT 163.420 10.460 165.720 10.700 ;
        RECT 163.420 10.350 163.870 10.460 ;
        RECT 165.270 10.350 165.720 10.460 ;
        RECT 166.670 10.700 167.120 10.800 ;
        RECT 168.520 10.700 168.970 10.800 ;
        RECT 166.670 10.460 168.970 10.700 ;
        RECT 166.670 10.380 167.120 10.460 ;
        RECT 147.180 9.800 148.710 10.010 ;
        RECT 149.090 9.800 149.540 9.890 ;
        RECT 149.920 9.800 151.450 10.010 ;
        RECT 160.680 10.010 161.130 10.290 ;
        RECT 164.500 10.010 164.950 10.290 ;
        RECT 167.720 10.020 168.130 10.460 ;
        RECT 168.520 10.350 168.970 10.460 ;
        RECT 170.160 10.700 170.610 10.800 ;
        RECT 172.010 10.700 172.460 10.800 ;
        RECT 170.160 10.460 172.460 10.700 ;
        RECT 170.160 10.350 170.610 10.460 ;
        RECT 171.000 10.020 171.410 10.460 ;
        RECT 172.010 10.380 172.460 10.460 ;
        RECT 173.410 10.700 173.860 10.770 ;
        RECT 174.460 10.700 174.870 11.130 ;
        RECT 175.260 10.700 175.710 10.800 ;
        RECT 173.410 10.460 175.710 10.700 ;
        RECT 173.410 10.350 173.860 10.460 ;
        RECT 175.260 10.350 175.710 10.460 ;
        RECT 176.920 10.700 177.370 10.800 ;
        RECT 177.760 10.700 178.170 11.130 ;
        RECT 180.920 11.060 182.470 11.280 ;
        RECT 182.850 11.270 183.280 11.330 ;
        RECT 183.660 11.280 184.110 11.330 ;
        RECT 184.710 11.280 185.210 11.670 ;
        RECT 183.660 11.060 185.210 11.280 ;
        RECT 194.420 11.670 195.970 11.890 ;
        RECT 194.420 11.280 194.920 11.670 ;
        RECT 195.520 11.620 195.970 11.670 ;
        RECT 196.350 11.620 196.780 11.680 ;
        RECT 197.160 11.670 198.710 11.890 ;
        RECT 201.460 11.820 201.870 12.250 ;
        RECT 202.260 12.150 202.710 12.250 ;
        RECT 203.920 12.490 204.370 12.600 ;
        RECT 205.770 12.490 206.220 12.600 ;
        RECT 203.920 12.250 206.220 12.490 ;
        RECT 203.920 12.150 204.370 12.250 ;
        RECT 204.760 11.820 205.170 12.250 ;
        RECT 205.770 12.180 206.220 12.250 ;
        RECT 207.170 12.490 207.620 12.570 ;
        RECT 208.220 12.490 208.630 12.930 ;
        RECT 209.020 12.490 209.470 12.600 ;
        RECT 207.170 12.250 209.470 12.490 ;
        RECT 207.170 12.150 207.620 12.250 ;
        RECT 209.020 12.150 209.470 12.250 ;
        RECT 210.660 12.490 211.110 12.600 ;
        RECT 211.500 12.490 211.910 12.930 ;
        RECT 214.680 12.660 215.130 12.940 ;
        RECT 212.510 12.490 212.960 12.570 ;
        RECT 210.660 12.250 212.960 12.490 ;
        RECT 210.660 12.150 211.110 12.250 ;
        RECT 212.510 12.150 212.960 12.250 ;
        RECT 213.910 12.490 214.360 12.600 ;
        RECT 215.760 12.490 216.210 12.600 ;
        RECT 213.910 12.250 216.210 12.490 ;
        RECT 213.910 12.180 214.360 12.250 ;
        RECT 197.160 11.620 197.610 11.670 ;
        RECT 195.520 11.330 197.610 11.620 ;
        RECT 195.520 11.280 195.970 11.330 ;
        RECT 178.770 10.700 179.220 10.770 ;
        RECT 176.920 10.460 179.220 10.700 ;
        RECT 176.920 10.350 177.370 10.460 ;
        RECT 178.770 10.350 179.220 10.460 ;
        RECT 180.170 10.700 180.620 10.800 ;
        RECT 182.020 10.700 182.470 10.800 ;
        RECT 180.170 10.460 182.470 10.700 ;
        RECT 180.170 10.380 180.620 10.460 ;
        RECT 160.680 9.800 162.210 10.010 ;
        RECT 162.590 9.800 163.040 9.890 ;
        RECT 163.420 9.800 164.950 10.010 ;
        RECT 174.180 10.010 174.630 10.290 ;
        RECT 178.000 10.010 178.450 10.290 ;
        RECT 181.220 10.020 181.630 10.460 ;
        RECT 182.020 10.350 182.470 10.460 ;
        RECT 183.660 10.700 184.110 10.800 ;
        RECT 185.510 10.700 185.960 10.800 ;
        RECT 183.660 10.460 185.960 10.700 ;
        RECT 183.660 10.350 184.110 10.460 ;
        RECT 184.500 10.020 184.910 10.460 ;
        RECT 185.510 10.380 185.960 10.460 ;
        RECT 186.910 10.700 187.360 10.770 ;
        RECT 187.960 10.700 188.370 11.130 ;
        RECT 188.760 10.700 189.210 10.800 ;
        RECT 186.910 10.460 189.210 10.700 ;
        RECT 186.910 10.350 187.360 10.460 ;
        RECT 188.760 10.350 189.210 10.460 ;
        RECT 190.420 10.700 190.870 10.800 ;
        RECT 191.260 10.700 191.670 11.130 ;
        RECT 194.420 11.060 195.970 11.280 ;
        RECT 196.350 11.270 196.780 11.330 ;
        RECT 197.160 11.280 197.610 11.330 ;
        RECT 198.210 11.280 198.710 11.670 ;
        RECT 197.160 11.060 198.710 11.280 ;
        RECT 207.920 11.670 209.470 11.890 ;
        RECT 207.920 11.280 208.420 11.670 ;
        RECT 209.020 11.620 209.470 11.670 ;
        RECT 209.850 11.620 210.280 11.680 ;
        RECT 210.660 11.670 212.210 11.890 ;
        RECT 214.960 11.820 215.370 12.250 ;
        RECT 215.760 12.150 216.210 12.250 ;
        RECT 210.660 11.620 211.110 11.670 ;
        RECT 209.020 11.330 211.110 11.620 ;
        RECT 209.020 11.280 209.470 11.330 ;
        RECT 192.270 10.700 192.720 10.770 ;
        RECT 190.420 10.460 192.720 10.700 ;
        RECT 190.420 10.350 190.870 10.460 ;
        RECT 192.270 10.350 192.720 10.460 ;
        RECT 193.670 10.700 194.120 10.800 ;
        RECT 195.520 10.700 195.970 10.800 ;
        RECT 193.670 10.460 195.970 10.700 ;
        RECT 193.670 10.380 194.120 10.460 ;
        RECT 174.180 9.800 175.710 10.010 ;
        RECT 176.090 9.800 176.540 9.890 ;
        RECT 176.920 9.800 178.450 10.010 ;
        RECT 187.680 10.010 188.130 10.290 ;
        RECT 191.500 10.010 191.950 10.290 ;
        RECT 194.720 10.020 195.130 10.460 ;
        RECT 195.520 10.350 195.970 10.460 ;
        RECT 197.160 10.700 197.610 10.800 ;
        RECT 199.010 10.700 199.460 10.800 ;
        RECT 197.160 10.460 199.460 10.700 ;
        RECT 197.160 10.350 197.610 10.460 ;
        RECT 198.000 10.020 198.410 10.460 ;
        RECT 199.010 10.380 199.460 10.460 ;
        RECT 200.410 10.700 200.860 10.770 ;
        RECT 201.460 10.700 201.870 11.130 ;
        RECT 202.260 10.700 202.710 10.800 ;
        RECT 200.410 10.460 202.710 10.700 ;
        RECT 200.410 10.350 200.860 10.460 ;
        RECT 202.260 10.350 202.710 10.460 ;
        RECT 203.920 10.700 204.370 10.800 ;
        RECT 204.760 10.700 205.170 11.130 ;
        RECT 207.920 11.060 209.470 11.280 ;
        RECT 209.850 11.270 210.280 11.330 ;
        RECT 210.660 11.280 211.110 11.330 ;
        RECT 211.710 11.280 212.210 11.670 ;
        RECT 210.660 11.060 212.210 11.280 ;
        RECT 205.770 10.700 206.220 10.770 ;
        RECT 203.920 10.460 206.220 10.700 ;
        RECT 203.920 10.350 204.370 10.460 ;
        RECT 205.770 10.350 206.220 10.460 ;
        RECT 207.170 10.700 207.620 10.800 ;
        RECT 209.020 10.700 209.470 10.800 ;
        RECT 207.170 10.460 209.470 10.700 ;
        RECT 207.170 10.380 207.620 10.460 ;
        RECT 187.680 9.800 189.210 10.010 ;
        RECT 189.590 9.800 190.040 9.890 ;
        RECT 190.420 9.800 191.950 10.010 ;
        RECT 201.180 10.010 201.630 10.290 ;
        RECT 205.000 10.010 205.450 10.290 ;
        RECT 208.220 10.020 208.630 10.460 ;
        RECT 209.020 10.350 209.470 10.460 ;
        RECT 210.660 10.700 211.110 10.800 ;
        RECT 212.510 10.700 212.960 10.800 ;
        RECT 210.660 10.460 212.960 10.700 ;
        RECT 210.660 10.350 211.110 10.460 ;
        RECT 211.500 10.020 211.910 10.460 ;
        RECT 212.510 10.380 212.960 10.460 ;
        RECT 213.910 10.700 214.360 10.770 ;
        RECT 214.960 10.700 215.370 11.130 ;
        RECT 215.760 10.700 216.210 10.800 ;
        RECT 213.910 10.460 216.210 10.700 ;
        RECT 213.910 10.350 214.360 10.460 ;
        RECT 215.760 10.350 216.210 10.460 ;
        RECT 201.180 9.800 202.710 10.010 ;
        RECT 203.090 9.800 203.540 9.890 ;
        RECT 203.920 9.800 205.450 10.010 ;
        RECT 214.680 10.010 215.130 10.290 ;
        RECT 214.680 9.800 216.210 10.010 ;
        RECT 216.590 9.800 217.030 9.890 ;
        RECT 13.260 9.540 15.370 9.800 ;
        RECT 26.760 9.540 28.870 9.800 ;
        RECT 40.260 9.540 42.370 9.800 ;
        RECT 53.760 9.540 55.870 9.800 ;
        RECT 67.260 9.540 69.370 9.800 ;
        RECT 80.760 9.540 82.870 9.800 ;
        RECT 94.260 9.540 96.370 9.800 ;
        RECT 107.760 9.540 109.870 9.800 ;
        RECT 121.260 9.540 123.370 9.800 ;
        RECT 134.760 9.540 136.870 9.800 ;
        RECT 148.260 9.540 150.370 9.800 ;
        RECT 161.760 9.540 163.870 9.800 ;
        RECT 175.260 9.540 177.370 9.800 ;
        RECT 188.760 9.540 190.870 9.800 ;
        RECT 202.260 9.540 204.370 9.800 ;
        RECT 215.760 9.540 217.030 9.800 ;
        RECT 12.180 9.330 13.710 9.540 ;
        RECT 14.090 9.450 14.540 9.540 ;
        RECT 14.920 9.330 16.450 9.540 ;
        RECT 1.420 8.880 1.870 8.990 ;
        RECT 3.270 8.880 3.720 8.990 ;
        RECT 1.420 8.640 3.720 8.880 ;
        RECT 1.420 8.540 1.870 8.640 ;
        RECT 2.260 8.210 2.670 8.640 ;
        RECT 3.270 8.570 3.720 8.640 ;
        RECT 4.670 8.880 5.120 8.960 ;
        RECT 5.720 8.880 6.130 9.320 ;
        RECT 6.520 8.880 6.970 8.990 ;
        RECT 4.670 8.640 6.970 8.880 ;
        RECT 4.670 8.540 5.120 8.640 ;
        RECT 6.520 8.540 6.970 8.640 ;
        RECT 8.160 8.880 8.610 8.990 ;
        RECT 9.000 8.880 9.410 9.320 ;
        RECT 12.180 9.050 12.630 9.330 ;
        RECT 16.000 9.050 16.450 9.330 ;
        RECT 25.680 9.330 27.210 9.540 ;
        RECT 27.590 9.450 28.040 9.540 ;
        RECT 28.420 9.330 29.950 9.540 ;
        RECT 10.010 8.880 10.460 8.960 ;
        RECT 8.160 8.640 10.460 8.880 ;
        RECT 8.160 8.540 8.610 8.640 ;
        RECT 10.010 8.540 10.460 8.640 ;
        RECT 11.410 8.880 11.860 8.990 ;
        RECT 13.260 8.880 13.710 8.990 ;
        RECT 11.410 8.640 13.710 8.880 ;
        RECT 11.410 8.570 11.860 8.640 ;
        RECT 5.420 8.060 6.970 8.280 ;
        RECT 5.420 7.670 5.920 8.060 ;
        RECT 6.520 8.010 6.970 8.060 ;
        RECT 7.350 8.010 7.780 8.070 ;
        RECT 8.160 8.060 9.710 8.280 ;
        RECT 12.460 8.210 12.870 8.640 ;
        RECT 13.260 8.540 13.710 8.640 ;
        RECT 14.920 8.880 15.370 8.990 ;
        RECT 16.770 8.880 17.220 8.990 ;
        RECT 14.920 8.640 17.220 8.880 ;
        RECT 14.920 8.540 15.370 8.640 ;
        RECT 15.760 8.210 16.170 8.640 ;
        RECT 16.770 8.570 17.220 8.640 ;
        RECT 18.170 8.880 18.620 8.960 ;
        RECT 19.220 8.880 19.630 9.320 ;
        RECT 20.020 8.880 20.470 8.990 ;
        RECT 18.170 8.640 20.470 8.880 ;
        RECT 18.170 8.540 18.620 8.640 ;
        RECT 20.020 8.540 20.470 8.640 ;
        RECT 21.660 8.880 22.110 8.990 ;
        RECT 22.500 8.880 22.910 9.320 ;
        RECT 25.680 9.050 26.130 9.330 ;
        RECT 29.500 9.050 29.950 9.330 ;
        RECT 39.180 9.330 40.710 9.540 ;
        RECT 41.090 9.450 41.540 9.540 ;
        RECT 41.920 9.330 43.450 9.540 ;
        RECT 23.510 8.880 23.960 8.960 ;
        RECT 21.660 8.640 23.960 8.880 ;
        RECT 21.660 8.540 22.110 8.640 ;
        RECT 23.510 8.540 23.960 8.640 ;
        RECT 24.910 8.880 25.360 8.990 ;
        RECT 26.760 8.880 27.210 8.990 ;
        RECT 24.910 8.640 27.210 8.880 ;
        RECT 24.910 8.570 25.360 8.640 ;
        RECT 8.160 8.010 8.610 8.060 ;
        RECT 6.520 7.720 8.610 8.010 ;
        RECT 6.520 7.670 6.970 7.720 ;
        RECT 1.420 7.090 1.870 7.190 ;
        RECT 2.260 7.090 2.670 7.520 ;
        RECT 5.420 7.450 6.970 7.670 ;
        RECT 7.350 7.660 7.780 7.720 ;
        RECT 8.160 7.670 8.610 7.720 ;
        RECT 9.210 7.670 9.710 8.060 ;
        RECT 8.160 7.450 9.710 7.670 ;
        RECT 18.920 8.060 20.470 8.280 ;
        RECT 18.920 7.670 19.420 8.060 ;
        RECT 20.020 8.010 20.470 8.060 ;
        RECT 20.850 8.010 21.280 8.070 ;
        RECT 21.660 8.060 23.210 8.280 ;
        RECT 25.960 8.210 26.370 8.640 ;
        RECT 26.760 8.540 27.210 8.640 ;
        RECT 28.420 8.880 28.870 8.990 ;
        RECT 30.270 8.880 30.720 8.990 ;
        RECT 28.420 8.640 30.720 8.880 ;
        RECT 28.420 8.540 28.870 8.640 ;
        RECT 29.260 8.210 29.670 8.640 ;
        RECT 30.270 8.570 30.720 8.640 ;
        RECT 31.670 8.880 32.120 8.960 ;
        RECT 32.720 8.880 33.130 9.320 ;
        RECT 33.520 8.880 33.970 8.990 ;
        RECT 31.670 8.640 33.970 8.880 ;
        RECT 31.670 8.540 32.120 8.640 ;
        RECT 33.520 8.540 33.970 8.640 ;
        RECT 35.160 8.880 35.610 8.990 ;
        RECT 36.000 8.880 36.410 9.320 ;
        RECT 39.180 9.050 39.630 9.330 ;
        RECT 43.000 9.050 43.450 9.330 ;
        RECT 52.680 9.330 54.210 9.540 ;
        RECT 54.590 9.450 55.040 9.540 ;
        RECT 55.420 9.330 56.950 9.540 ;
        RECT 37.010 8.880 37.460 8.960 ;
        RECT 35.160 8.640 37.460 8.880 ;
        RECT 35.160 8.540 35.610 8.640 ;
        RECT 37.010 8.540 37.460 8.640 ;
        RECT 38.410 8.880 38.860 8.990 ;
        RECT 40.260 8.880 40.710 8.990 ;
        RECT 38.410 8.640 40.710 8.880 ;
        RECT 38.410 8.570 38.860 8.640 ;
        RECT 21.660 8.010 22.110 8.060 ;
        RECT 20.020 7.720 22.110 8.010 ;
        RECT 20.020 7.670 20.470 7.720 ;
        RECT 3.270 7.090 3.720 7.160 ;
        RECT 1.420 6.850 3.720 7.090 ;
        RECT 1.420 6.740 1.870 6.850 ;
        RECT 3.270 6.740 3.720 6.850 ;
        RECT 4.670 7.090 5.120 7.190 ;
        RECT 6.520 7.090 6.970 7.190 ;
        RECT 4.670 6.850 6.970 7.090 ;
        RECT 4.670 6.770 5.120 6.850 ;
        RECT 5.720 6.410 6.130 6.850 ;
        RECT 6.520 6.740 6.970 6.850 ;
        RECT 8.160 7.090 8.610 7.190 ;
        RECT 10.010 7.090 10.460 7.190 ;
        RECT 8.160 6.850 10.460 7.090 ;
        RECT 8.160 6.740 8.610 6.850 ;
        RECT 9.000 6.410 9.410 6.850 ;
        RECT 10.010 6.770 10.460 6.850 ;
        RECT 11.410 7.090 11.860 7.160 ;
        RECT 12.460 7.090 12.870 7.520 ;
        RECT 13.260 7.090 13.710 7.190 ;
        RECT 11.410 6.850 13.710 7.090 ;
        RECT 11.410 6.740 11.860 6.850 ;
        RECT 13.260 6.740 13.710 6.850 ;
        RECT 14.920 7.090 15.370 7.190 ;
        RECT 15.760 7.090 16.170 7.520 ;
        RECT 18.920 7.450 20.470 7.670 ;
        RECT 20.850 7.660 21.280 7.720 ;
        RECT 21.660 7.670 22.110 7.720 ;
        RECT 22.710 7.670 23.210 8.060 ;
        RECT 21.660 7.450 23.210 7.670 ;
        RECT 32.420 8.060 33.970 8.280 ;
        RECT 32.420 7.670 32.920 8.060 ;
        RECT 33.520 8.010 33.970 8.060 ;
        RECT 34.350 8.010 34.780 8.070 ;
        RECT 35.160 8.060 36.710 8.280 ;
        RECT 39.460 8.210 39.870 8.640 ;
        RECT 40.260 8.540 40.710 8.640 ;
        RECT 41.920 8.880 42.370 8.990 ;
        RECT 43.770 8.880 44.220 8.990 ;
        RECT 41.920 8.640 44.220 8.880 ;
        RECT 41.920 8.540 42.370 8.640 ;
        RECT 42.760 8.210 43.170 8.640 ;
        RECT 43.770 8.570 44.220 8.640 ;
        RECT 45.170 8.880 45.620 8.960 ;
        RECT 46.220 8.880 46.630 9.320 ;
        RECT 47.020 8.880 47.470 8.990 ;
        RECT 45.170 8.640 47.470 8.880 ;
        RECT 45.170 8.540 45.620 8.640 ;
        RECT 47.020 8.540 47.470 8.640 ;
        RECT 48.660 8.880 49.110 8.990 ;
        RECT 49.500 8.880 49.910 9.320 ;
        RECT 52.680 9.050 53.130 9.330 ;
        RECT 56.500 9.050 56.950 9.330 ;
        RECT 66.180 9.330 67.710 9.540 ;
        RECT 68.090 9.450 68.540 9.540 ;
        RECT 68.920 9.330 70.450 9.540 ;
        RECT 50.510 8.880 50.960 8.960 ;
        RECT 48.660 8.640 50.960 8.880 ;
        RECT 48.660 8.540 49.110 8.640 ;
        RECT 50.510 8.540 50.960 8.640 ;
        RECT 51.910 8.880 52.360 8.990 ;
        RECT 53.760 8.880 54.210 8.990 ;
        RECT 51.910 8.640 54.210 8.880 ;
        RECT 51.910 8.570 52.360 8.640 ;
        RECT 35.160 8.010 35.610 8.060 ;
        RECT 33.520 7.720 35.610 8.010 ;
        RECT 33.520 7.670 33.970 7.720 ;
        RECT 16.770 7.090 17.220 7.160 ;
        RECT 14.920 6.850 17.220 7.090 ;
        RECT 14.920 6.740 15.370 6.850 ;
        RECT 16.770 6.740 17.220 6.850 ;
        RECT 18.170 7.090 18.620 7.190 ;
        RECT 20.020 7.090 20.470 7.190 ;
        RECT 18.170 6.850 20.470 7.090 ;
        RECT 18.170 6.770 18.620 6.850 ;
        RECT 12.180 6.400 12.630 6.680 ;
        RECT 16.000 6.400 16.450 6.680 ;
        RECT 19.220 6.410 19.630 6.850 ;
        RECT 20.020 6.740 20.470 6.850 ;
        RECT 21.660 7.090 22.110 7.190 ;
        RECT 23.510 7.090 23.960 7.190 ;
        RECT 21.660 6.850 23.960 7.090 ;
        RECT 21.660 6.740 22.110 6.850 ;
        RECT 22.500 6.410 22.910 6.850 ;
        RECT 23.510 6.770 23.960 6.850 ;
        RECT 24.910 7.090 25.360 7.160 ;
        RECT 25.960 7.090 26.370 7.520 ;
        RECT 26.760 7.090 27.210 7.190 ;
        RECT 24.910 6.850 27.210 7.090 ;
        RECT 24.910 6.740 25.360 6.850 ;
        RECT 26.760 6.740 27.210 6.850 ;
        RECT 28.420 7.090 28.870 7.190 ;
        RECT 29.260 7.090 29.670 7.520 ;
        RECT 32.420 7.450 33.970 7.670 ;
        RECT 34.350 7.660 34.780 7.720 ;
        RECT 35.160 7.670 35.610 7.720 ;
        RECT 36.210 7.670 36.710 8.060 ;
        RECT 35.160 7.450 36.710 7.670 ;
        RECT 45.920 8.060 47.470 8.280 ;
        RECT 45.920 7.670 46.420 8.060 ;
        RECT 47.020 8.010 47.470 8.060 ;
        RECT 47.850 8.010 48.280 8.070 ;
        RECT 48.660 8.060 50.210 8.280 ;
        RECT 52.960 8.210 53.370 8.640 ;
        RECT 53.760 8.540 54.210 8.640 ;
        RECT 55.420 8.880 55.870 8.990 ;
        RECT 57.270 8.880 57.720 8.990 ;
        RECT 55.420 8.640 57.720 8.880 ;
        RECT 55.420 8.540 55.870 8.640 ;
        RECT 56.260 8.210 56.670 8.640 ;
        RECT 57.270 8.570 57.720 8.640 ;
        RECT 58.670 8.880 59.120 8.960 ;
        RECT 59.720 8.880 60.130 9.320 ;
        RECT 60.520 8.880 60.970 8.990 ;
        RECT 58.670 8.640 60.970 8.880 ;
        RECT 58.670 8.540 59.120 8.640 ;
        RECT 60.520 8.540 60.970 8.640 ;
        RECT 62.160 8.880 62.610 8.990 ;
        RECT 63.000 8.880 63.410 9.320 ;
        RECT 66.180 9.050 66.630 9.330 ;
        RECT 70.000 9.050 70.450 9.330 ;
        RECT 79.680 9.330 81.210 9.540 ;
        RECT 81.590 9.450 82.040 9.540 ;
        RECT 82.420 9.330 83.950 9.540 ;
        RECT 64.010 8.880 64.460 8.960 ;
        RECT 62.160 8.640 64.460 8.880 ;
        RECT 62.160 8.540 62.610 8.640 ;
        RECT 64.010 8.540 64.460 8.640 ;
        RECT 65.410 8.880 65.860 8.990 ;
        RECT 67.260 8.880 67.710 8.990 ;
        RECT 65.410 8.640 67.710 8.880 ;
        RECT 65.410 8.570 65.860 8.640 ;
        RECT 48.660 8.010 49.110 8.060 ;
        RECT 47.020 7.720 49.110 8.010 ;
        RECT 47.020 7.670 47.470 7.720 ;
        RECT 30.270 7.090 30.720 7.160 ;
        RECT 28.420 6.850 30.720 7.090 ;
        RECT 28.420 6.740 28.870 6.850 ;
        RECT 30.270 6.740 30.720 6.850 ;
        RECT 31.670 7.090 32.120 7.190 ;
        RECT 33.520 7.090 33.970 7.190 ;
        RECT 31.670 6.850 33.970 7.090 ;
        RECT 31.670 6.770 32.120 6.850 ;
        RECT 12.180 6.190 13.710 6.400 ;
        RECT 14.090 6.190 14.540 6.280 ;
        RECT 14.920 6.190 16.450 6.400 ;
        RECT 25.680 6.400 26.130 6.680 ;
        RECT 29.500 6.400 29.950 6.680 ;
        RECT 32.720 6.410 33.130 6.850 ;
        RECT 33.520 6.740 33.970 6.850 ;
        RECT 35.160 7.090 35.610 7.190 ;
        RECT 37.010 7.090 37.460 7.190 ;
        RECT 35.160 6.850 37.460 7.090 ;
        RECT 35.160 6.740 35.610 6.850 ;
        RECT 36.000 6.410 36.410 6.850 ;
        RECT 37.010 6.770 37.460 6.850 ;
        RECT 38.410 7.090 38.860 7.160 ;
        RECT 39.460 7.090 39.870 7.520 ;
        RECT 40.260 7.090 40.710 7.190 ;
        RECT 38.410 6.850 40.710 7.090 ;
        RECT 38.410 6.740 38.860 6.850 ;
        RECT 40.260 6.740 40.710 6.850 ;
        RECT 41.920 7.090 42.370 7.190 ;
        RECT 42.760 7.090 43.170 7.520 ;
        RECT 45.920 7.450 47.470 7.670 ;
        RECT 47.850 7.660 48.280 7.720 ;
        RECT 48.660 7.670 49.110 7.720 ;
        RECT 49.710 7.670 50.210 8.060 ;
        RECT 48.660 7.450 50.210 7.670 ;
        RECT 59.420 8.060 60.970 8.280 ;
        RECT 59.420 7.670 59.920 8.060 ;
        RECT 60.520 8.010 60.970 8.060 ;
        RECT 61.350 8.010 61.780 8.070 ;
        RECT 62.160 8.060 63.710 8.280 ;
        RECT 66.460 8.210 66.870 8.640 ;
        RECT 67.260 8.540 67.710 8.640 ;
        RECT 68.920 8.880 69.370 8.990 ;
        RECT 70.770 8.880 71.220 8.990 ;
        RECT 68.920 8.640 71.220 8.880 ;
        RECT 68.920 8.540 69.370 8.640 ;
        RECT 69.760 8.210 70.170 8.640 ;
        RECT 70.770 8.570 71.220 8.640 ;
        RECT 72.170 8.880 72.620 8.960 ;
        RECT 73.220 8.880 73.630 9.320 ;
        RECT 74.020 8.880 74.470 8.990 ;
        RECT 72.170 8.640 74.470 8.880 ;
        RECT 72.170 8.540 72.620 8.640 ;
        RECT 74.020 8.540 74.470 8.640 ;
        RECT 75.660 8.880 76.110 8.990 ;
        RECT 76.500 8.880 76.910 9.320 ;
        RECT 79.680 9.050 80.130 9.330 ;
        RECT 83.500 9.050 83.950 9.330 ;
        RECT 93.180 9.330 94.710 9.540 ;
        RECT 95.090 9.450 95.540 9.540 ;
        RECT 95.920 9.330 97.450 9.540 ;
        RECT 77.510 8.880 77.960 8.960 ;
        RECT 75.660 8.640 77.960 8.880 ;
        RECT 75.660 8.540 76.110 8.640 ;
        RECT 77.510 8.540 77.960 8.640 ;
        RECT 78.910 8.880 79.360 8.990 ;
        RECT 80.760 8.880 81.210 8.990 ;
        RECT 78.910 8.640 81.210 8.880 ;
        RECT 78.910 8.570 79.360 8.640 ;
        RECT 62.160 8.010 62.610 8.060 ;
        RECT 60.520 7.720 62.610 8.010 ;
        RECT 60.520 7.670 60.970 7.720 ;
        RECT 43.770 7.090 44.220 7.160 ;
        RECT 41.920 6.850 44.220 7.090 ;
        RECT 41.920 6.740 42.370 6.850 ;
        RECT 43.770 6.740 44.220 6.850 ;
        RECT 45.170 7.090 45.620 7.190 ;
        RECT 47.020 7.090 47.470 7.190 ;
        RECT 45.170 6.850 47.470 7.090 ;
        RECT 45.170 6.770 45.620 6.850 ;
        RECT 25.680 6.190 27.210 6.400 ;
        RECT 27.590 6.190 28.040 6.280 ;
        RECT 28.420 6.190 29.950 6.400 ;
        RECT 39.180 6.400 39.630 6.680 ;
        RECT 43.000 6.400 43.450 6.680 ;
        RECT 46.220 6.410 46.630 6.850 ;
        RECT 47.020 6.740 47.470 6.850 ;
        RECT 48.660 7.090 49.110 7.190 ;
        RECT 50.510 7.090 50.960 7.190 ;
        RECT 48.660 6.850 50.960 7.090 ;
        RECT 48.660 6.740 49.110 6.850 ;
        RECT 49.500 6.410 49.910 6.850 ;
        RECT 50.510 6.770 50.960 6.850 ;
        RECT 51.910 7.090 52.360 7.160 ;
        RECT 52.960 7.090 53.370 7.520 ;
        RECT 53.760 7.090 54.210 7.190 ;
        RECT 51.910 6.850 54.210 7.090 ;
        RECT 51.910 6.740 52.360 6.850 ;
        RECT 53.760 6.740 54.210 6.850 ;
        RECT 55.420 7.090 55.870 7.190 ;
        RECT 56.260 7.090 56.670 7.520 ;
        RECT 59.420 7.450 60.970 7.670 ;
        RECT 61.350 7.660 61.780 7.720 ;
        RECT 62.160 7.670 62.610 7.720 ;
        RECT 63.210 7.670 63.710 8.060 ;
        RECT 62.160 7.450 63.710 7.670 ;
        RECT 72.920 8.060 74.470 8.280 ;
        RECT 72.920 7.670 73.420 8.060 ;
        RECT 74.020 8.010 74.470 8.060 ;
        RECT 74.850 8.010 75.280 8.070 ;
        RECT 75.660 8.060 77.210 8.280 ;
        RECT 79.960 8.210 80.370 8.640 ;
        RECT 80.760 8.540 81.210 8.640 ;
        RECT 82.420 8.880 82.870 8.990 ;
        RECT 84.270 8.880 84.720 8.990 ;
        RECT 82.420 8.640 84.720 8.880 ;
        RECT 82.420 8.540 82.870 8.640 ;
        RECT 83.260 8.210 83.670 8.640 ;
        RECT 84.270 8.570 84.720 8.640 ;
        RECT 85.670 8.880 86.120 8.960 ;
        RECT 86.720 8.880 87.130 9.320 ;
        RECT 87.520 8.880 87.970 8.990 ;
        RECT 85.670 8.640 87.970 8.880 ;
        RECT 85.670 8.540 86.120 8.640 ;
        RECT 87.520 8.540 87.970 8.640 ;
        RECT 89.160 8.880 89.610 8.990 ;
        RECT 90.000 8.880 90.410 9.320 ;
        RECT 93.180 9.050 93.630 9.330 ;
        RECT 97.000 9.050 97.450 9.330 ;
        RECT 106.680 9.330 108.210 9.540 ;
        RECT 108.590 9.450 109.040 9.540 ;
        RECT 109.420 9.330 110.950 9.540 ;
        RECT 91.010 8.880 91.460 8.960 ;
        RECT 89.160 8.640 91.460 8.880 ;
        RECT 89.160 8.540 89.610 8.640 ;
        RECT 91.010 8.540 91.460 8.640 ;
        RECT 92.410 8.880 92.860 8.990 ;
        RECT 94.260 8.880 94.710 8.990 ;
        RECT 92.410 8.640 94.710 8.880 ;
        RECT 92.410 8.570 92.860 8.640 ;
        RECT 75.660 8.010 76.110 8.060 ;
        RECT 74.020 7.720 76.110 8.010 ;
        RECT 74.020 7.670 74.470 7.720 ;
        RECT 57.270 7.090 57.720 7.160 ;
        RECT 55.420 6.850 57.720 7.090 ;
        RECT 55.420 6.740 55.870 6.850 ;
        RECT 57.270 6.740 57.720 6.850 ;
        RECT 58.670 7.090 59.120 7.190 ;
        RECT 60.520 7.090 60.970 7.190 ;
        RECT 58.670 6.850 60.970 7.090 ;
        RECT 58.670 6.770 59.120 6.850 ;
        RECT 39.180 6.190 40.710 6.400 ;
        RECT 41.090 6.190 41.540 6.280 ;
        RECT 41.920 6.190 43.450 6.400 ;
        RECT 52.680 6.400 53.130 6.680 ;
        RECT 56.500 6.400 56.950 6.680 ;
        RECT 59.720 6.410 60.130 6.850 ;
        RECT 60.520 6.740 60.970 6.850 ;
        RECT 62.160 7.090 62.610 7.190 ;
        RECT 64.010 7.090 64.460 7.190 ;
        RECT 62.160 6.850 64.460 7.090 ;
        RECT 62.160 6.740 62.610 6.850 ;
        RECT 63.000 6.410 63.410 6.850 ;
        RECT 64.010 6.770 64.460 6.850 ;
        RECT 65.410 7.090 65.860 7.160 ;
        RECT 66.460 7.090 66.870 7.520 ;
        RECT 67.260 7.090 67.710 7.190 ;
        RECT 65.410 6.850 67.710 7.090 ;
        RECT 65.410 6.740 65.860 6.850 ;
        RECT 67.260 6.740 67.710 6.850 ;
        RECT 68.920 7.090 69.370 7.190 ;
        RECT 69.760 7.090 70.170 7.520 ;
        RECT 72.920 7.450 74.470 7.670 ;
        RECT 74.850 7.660 75.280 7.720 ;
        RECT 75.660 7.670 76.110 7.720 ;
        RECT 76.710 7.670 77.210 8.060 ;
        RECT 75.660 7.450 77.210 7.670 ;
        RECT 86.420 8.060 87.970 8.280 ;
        RECT 86.420 7.670 86.920 8.060 ;
        RECT 87.520 8.010 87.970 8.060 ;
        RECT 88.350 8.010 88.780 8.070 ;
        RECT 89.160 8.060 90.710 8.280 ;
        RECT 93.460 8.210 93.870 8.640 ;
        RECT 94.260 8.540 94.710 8.640 ;
        RECT 95.920 8.880 96.370 8.990 ;
        RECT 97.770 8.880 98.220 8.990 ;
        RECT 95.920 8.640 98.220 8.880 ;
        RECT 95.920 8.540 96.370 8.640 ;
        RECT 96.760 8.210 97.170 8.640 ;
        RECT 97.770 8.570 98.220 8.640 ;
        RECT 99.170 8.880 99.620 8.960 ;
        RECT 100.220 8.880 100.630 9.320 ;
        RECT 101.020 8.880 101.470 8.990 ;
        RECT 99.170 8.640 101.470 8.880 ;
        RECT 99.170 8.540 99.620 8.640 ;
        RECT 101.020 8.540 101.470 8.640 ;
        RECT 102.660 8.880 103.110 8.990 ;
        RECT 103.500 8.880 103.910 9.320 ;
        RECT 106.680 9.050 107.130 9.330 ;
        RECT 110.500 9.050 110.950 9.330 ;
        RECT 120.180 9.330 121.710 9.540 ;
        RECT 122.090 9.450 122.540 9.540 ;
        RECT 122.920 9.330 124.450 9.540 ;
        RECT 104.510 8.880 104.960 8.960 ;
        RECT 102.660 8.640 104.960 8.880 ;
        RECT 102.660 8.540 103.110 8.640 ;
        RECT 104.510 8.540 104.960 8.640 ;
        RECT 105.910 8.880 106.360 8.990 ;
        RECT 107.760 8.880 108.210 8.990 ;
        RECT 105.910 8.640 108.210 8.880 ;
        RECT 105.910 8.570 106.360 8.640 ;
        RECT 89.160 8.010 89.610 8.060 ;
        RECT 87.520 7.720 89.610 8.010 ;
        RECT 87.520 7.670 87.970 7.720 ;
        RECT 70.770 7.090 71.220 7.160 ;
        RECT 68.920 6.850 71.220 7.090 ;
        RECT 68.920 6.740 69.370 6.850 ;
        RECT 70.770 6.740 71.220 6.850 ;
        RECT 72.170 7.090 72.620 7.190 ;
        RECT 74.020 7.090 74.470 7.190 ;
        RECT 72.170 6.850 74.470 7.090 ;
        RECT 72.170 6.770 72.620 6.850 ;
        RECT 52.680 6.190 54.210 6.400 ;
        RECT 54.590 6.190 55.040 6.280 ;
        RECT 55.420 6.190 56.950 6.400 ;
        RECT 66.180 6.400 66.630 6.680 ;
        RECT 70.000 6.400 70.450 6.680 ;
        RECT 73.220 6.410 73.630 6.850 ;
        RECT 74.020 6.740 74.470 6.850 ;
        RECT 75.660 7.090 76.110 7.190 ;
        RECT 77.510 7.090 77.960 7.190 ;
        RECT 75.660 6.850 77.960 7.090 ;
        RECT 75.660 6.740 76.110 6.850 ;
        RECT 76.500 6.410 76.910 6.850 ;
        RECT 77.510 6.770 77.960 6.850 ;
        RECT 78.910 7.090 79.360 7.160 ;
        RECT 79.960 7.090 80.370 7.520 ;
        RECT 80.760 7.090 81.210 7.190 ;
        RECT 78.910 6.850 81.210 7.090 ;
        RECT 78.910 6.740 79.360 6.850 ;
        RECT 80.760 6.740 81.210 6.850 ;
        RECT 82.420 7.090 82.870 7.190 ;
        RECT 83.260 7.090 83.670 7.520 ;
        RECT 86.420 7.450 87.970 7.670 ;
        RECT 88.350 7.660 88.780 7.720 ;
        RECT 89.160 7.670 89.610 7.720 ;
        RECT 90.210 7.670 90.710 8.060 ;
        RECT 89.160 7.450 90.710 7.670 ;
        RECT 99.920 8.060 101.470 8.280 ;
        RECT 99.920 7.670 100.420 8.060 ;
        RECT 101.020 8.010 101.470 8.060 ;
        RECT 101.850 8.010 102.280 8.070 ;
        RECT 102.660 8.060 104.210 8.280 ;
        RECT 106.960 8.210 107.370 8.640 ;
        RECT 107.760 8.540 108.210 8.640 ;
        RECT 109.420 8.880 109.870 8.990 ;
        RECT 111.270 8.880 111.720 8.990 ;
        RECT 109.420 8.640 111.720 8.880 ;
        RECT 109.420 8.540 109.870 8.640 ;
        RECT 110.260 8.210 110.670 8.640 ;
        RECT 111.270 8.570 111.720 8.640 ;
        RECT 112.670 8.880 113.120 8.960 ;
        RECT 113.720 8.880 114.130 9.320 ;
        RECT 114.520 8.880 114.970 8.990 ;
        RECT 112.670 8.640 114.970 8.880 ;
        RECT 112.670 8.540 113.120 8.640 ;
        RECT 114.520 8.540 114.970 8.640 ;
        RECT 116.160 8.880 116.610 8.990 ;
        RECT 117.000 8.880 117.410 9.320 ;
        RECT 120.180 9.050 120.630 9.330 ;
        RECT 124.000 9.050 124.450 9.330 ;
        RECT 133.680 9.330 135.210 9.540 ;
        RECT 135.590 9.450 136.040 9.540 ;
        RECT 136.420 9.330 137.950 9.540 ;
        RECT 118.010 8.880 118.460 8.960 ;
        RECT 116.160 8.640 118.460 8.880 ;
        RECT 116.160 8.540 116.610 8.640 ;
        RECT 118.010 8.540 118.460 8.640 ;
        RECT 119.410 8.880 119.860 8.990 ;
        RECT 121.260 8.880 121.710 8.990 ;
        RECT 119.410 8.640 121.710 8.880 ;
        RECT 119.410 8.570 119.860 8.640 ;
        RECT 102.660 8.010 103.110 8.060 ;
        RECT 101.020 7.720 103.110 8.010 ;
        RECT 101.020 7.670 101.470 7.720 ;
        RECT 84.270 7.090 84.720 7.160 ;
        RECT 82.420 6.850 84.720 7.090 ;
        RECT 82.420 6.740 82.870 6.850 ;
        RECT 84.270 6.740 84.720 6.850 ;
        RECT 85.670 7.090 86.120 7.190 ;
        RECT 87.520 7.090 87.970 7.190 ;
        RECT 85.670 6.850 87.970 7.090 ;
        RECT 85.670 6.770 86.120 6.850 ;
        RECT 66.180 6.190 67.710 6.400 ;
        RECT 68.090 6.190 68.540 6.280 ;
        RECT 68.920 6.190 70.450 6.400 ;
        RECT 79.680 6.400 80.130 6.680 ;
        RECT 83.500 6.400 83.950 6.680 ;
        RECT 86.720 6.410 87.130 6.850 ;
        RECT 87.520 6.740 87.970 6.850 ;
        RECT 89.160 7.090 89.610 7.190 ;
        RECT 91.010 7.090 91.460 7.190 ;
        RECT 89.160 6.850 91.460 7.090 ;
        RECT 89.160 6.740 89.610 6.850 ;
        RECT 90.000 6.410 90.410 6.850 ;
        RECT 91.010 6.770 91.460 6.850 ;
        RECT 92.410 7.090 92.860 7.160 ;
        RECT 93.460 7.090 93.870 7.520 ;
        RECT 94.260 7.090 94.710 7.190 ;
        RECT 92.410 6.850 94.710 7.090 ;
        RECT 92.410 6.740 92.860 6.850 ;
        RECT 94.260 6.740 94.710 6.850 ;
        RECT 95.920 7.090 96.370 7.190 ;
        RECT 96.760 7.090 97.170 7.520 ;
        RECT 99.920 7.450 101.470 7.670 ;
        RECT 101.850 7.660 102.280 7.720 ;
        RECT 102.660 7.670 103.110 7.720 ;
        RECT 103.710 7.670 104.210 8.060 ;
        RECT 102.660 7.450 104.210 7.670 ;
        RECT 113.420 8.060 114.970 8.280 ;
        RECT 113.420 7.670 113.920 8.060 ;
        RECT 114.520 8.010 114.970 8.060 ;
        RECT 115.350 8.010 115.780 8.070 ;
        RECT 116.160 8.060 117.710 8.280 ;
        RECT 120.460 8.210 120.870 8.640 ;
        RECT 121.260 8.540 121.710 8.640 ;
        RECT 122.920 8.880 123.370 8.990 ;
        RECT 124.770 8.880 125.220 8.990 ;
        RECT 122.920 8.640 125.220 8.880 ;
        RECT 122.920 8.540 123.370 8.640 ;
        RECT 123.760 8.210 124.170 8.640 ;
        RECT 124.770 8.570 125.220 8.640 ;
        RECT 126.170 8.880 126.620 8.960 ;
        RECT 127.220 8.880 127.630 9.320 ;
        RECT 128.020 8.880 128.470 8.990 ;
        RECT 126.170 8.640 128.470 8.880 ;
        RECT 126.170 8.540 126.620 8.640 ;
        RECT 128.020 8.540 128.470 8.640 ;
        RECT 129.660 8.880 130.110 8.990 ;
        RECT 130.500 8.880 130.910 9.320 ;
        RECT 133.680 9.050 134.130 9.330 ;
        RECT 137.500 9.050 137.950 9.330 ;
        RECT 147.180 9.330 148.710 9.540 ;
        RECT 149.090 9.450 149.540 9.540 ;
        RECT 149.920 9.330 151.450 9.540 ;
        RECT 131.510 8.880 131.960 8.960 ;
        RECT 129.660 8.640 131.960 8.880 ;
        RECT 129.660 8.540 130.110 8.640 ;
        RECT 131.510 8.540 131.960 8.640 ;
        RECT 132.910 8.880 133.360 8.990 ;
        RECT 134.760 8.880 135.210 8.990 ;
        RECT 132.910 8.640 135.210 8.880 ;
        RECT 132.910 8.570 133.360 8.640 ;
        RECT 116.160 8.010 116.610 8.060 ;
        RECT 114.520 7.720 116.610 8.010 ;
        RECT 114.520 7.670 114.970 7.720 ;
        RECT 97.770 7.090 98.220 7.160 ;
        RECT 95.920 6.850 98.220 7.090 ;
        RECT 95.920 6.740 96.370 6.850 ;
        RECT 97.770 6.740 98.220 6.850 ;
        RECT 99.170 7.090 99.620 7.190 ;
        RECT 101.020 7.090 101.470 7.190 ;
        RECT 99.170 6.850 101.470 7.090 ;
        RECT 99.170 6.770 99.620 6.850 ;
        RECT 79.680 6.190 81.210 6.400 ;
        RECT 81.590 6.190 82.040 6.280 ;
        RECT 82.420 6.190 83.950 6.400 ;
        RECT 93.180 6.400 93.630 6.680 ;
        RECT 97.000 6.400 97.450 6.680 ;
        RECT 100.220 6.410 100.630 6.850 ;
        RECT 101.020 6.740 101.470 6.850 ;
        RECT 102.660 7.090 103.110 7.190 ;
        RECT 104.510 7.090 104.960 7.190 ;
        RECT 102.660 6.850 104.960 7.090 ;
        RECT 102.660 6.740 103.110 6.850 ;
        RECT 103.500 6.410 103.910 6.850 ;
        RECT 104.510 6.770 104.960 6.850 ;
        RECT 105.910 7.090 106.360 7.160 ;
        RECT 106.960 7.090 107.370 7.520 ;
        RECT 107.760 7.090 108.210 7.190 ;
        RECT 105.910 6.850 108.210 7.090 ;
        RECT 105.910 6.740 106.360 6.850 ;
        RECT 107.760 6.740 108.210 6.850 ;
        RECT 109.420 7.090 109.870 7.190 ;
        RECT 110.260 7.090 110.670 7.520 ;
        RECT 113.420 7.450 114.970 7.670 ;
        RECT 115.350 7.660 115.780 7.720 ;
        RECT 116.160 7.670 116.610 7.720 ;
        RECT 117.210 7.670 117.710 8.060 ;
        RECT 116.160 7.450 117.710 7.670 ;
        RECT 126.920 8.060 128.470 8.280 ;
        RECT 126.920 7.670 127.420 8.060 ;
        RECT 128.020 8.010 128.470 8.060 ;
        RECT 128.850 8.010 129.280 8.070 ;
        RECT 129.660 8.060 131.210 8.280 ;
        RECT 133.960 8.210 134.370 8.640 ;
        RECT 134.760 8.540 135.210 8.640 ;
        RECT 136.420 8.880 136.870 8.990 ;
        RECT 138.270 8.880 138.720 8.990 ;
        RECT 136.420 8.640 138.720 8.880 ;
        RECT 136.420 8.540 136.870 8.640 ;
        RECT 137.260 8.210 137.670 8.640 ;
        RECT 138.270 8.570 138.720 8.640 ;
        RECT 139.670 8.880 140.120 8.960 ;
        RECT 140.720 8.880 141.130 9.320 ;
        RECT 141.520 8.880 141.970 8.990 ;
        RECT 139.670 8.640 141.970 8.880 ;
        RECT 139.670 8.540 140.120 8.640 ;
        RECT 141.520 8.540 141.970 8.640 ;
        RECT 143.160 8.880 143.610 8.990 ;
        RECT 144.000 8.880 144.410 9.320 ;
        RECT 147.180 9.050 147.630 9.330 ;
        RECT 151.000 9.050 151.450 9.330 ;
        RECT 160.680 9.330 162.210 9.540 ;
        RECT 162.590 9.450 163.040 9.540 ;
        RECT 163.420 9.330 164.950 9.540 ;
        RECT 145.010 8.880 145.460 8.960 ;
        RECT 143.160 8.640 145.460 8.880 ;
        RECT 143.160 8.540 143.610 8.640 ;
        RECT 145.010 8.540 145.460 8.640 ;
        RECT 146.410 8.880 146.860 8.990 ;
        RECT 148.260 8.880 148.710 8.990 ;
        RECT 146.410 8.640 148.710 8.880 ;
        RECT 146.410 8.570 146.860 8.640 ;
        RECT 129.660 8.010 130.110 8.060 ;
        RECT 128.020 7.720 130.110 8.010 ;
        RECT 128.020 7.670 128.470 7.720 ;
        RECT 111.270 7.090 111.720 7.160 ;
        RECT 109.420 6.850 111.720 7.090 ;
        RECT 109.420 6.740 109.870 6.850 ;
        RECT 111.270 6.740 111.720 6.850 ;
        RECT 112.670 7.090 113.120 7.190 ;
        RECT 114.520 7.090 114.970 7.190 ;
        RECT 112.670 6.850 114.970 7.090 ;
        RECT 112.670 6.770 113.120 6.850 ;
        RECT 93.180 6.190 94.710 6.400 ;
        RECT 95.090 6.190 95.540 6.280 ;
        RECT 95.920 6.190 97.450 6.400 ;
        RECT 106.680 6.400 107.130 6.680 ;
        RECT 110.500 6.400 110.950 6.680 ;
        RECT 113.720 6.410 114.130 6.850 ;
        RECT 114.520 6.740 114.970 6.850 ;
        RECT 116.160 7.090 116.610 7.190 ;
        RECT 118.010 7.090 118.460 7.190 ;
        RECT 116.160 6.850 118.460 7.090 ;
        RECT 116.160 6.740 116.610 6.850 ;
        RECT 117.000 6.410 117.410 6.850 ;
        RECT 118.010 6.770 118.460 6.850 ;
        RECT 119.410 7.090 119.860 7.160 ;
        RECT 120.460 7.090 120.870 7.520 ;
        RECT 121.260 7.090 121.710 7.190 ;
        RECT 119.410 6.850 121.710 7.090 ;
        RECT 119.410 6.740 119.860 6.850 ;
        RECT 121.260 6.740 121.710 6.850 ;
        RECT 122.920 7.090 123.370 7.190 ;
        RECT 123.760 7.090 124.170 7.520 ;
        RECT 126.920 7.450 128.470 7.670 ;
        RECT 128.850 7.660 129.280 7.720 ;
        RECT 129.660 7.670 130.110 7.720 ;
        RECT 130.710 7.670 131.210 8.060 ;
        RECT 129.660 7.450 131.210 7.670 ;
        RECT 140.420 8.060 141.970 8.280 ;
        RECT 140.420 7.670 140.920 8.060 ;
        RECT 141.520 8.010 141.970 8.060 ;
        RECT 142.350 8.010 142.780 8.070 ;
        RECT 143.160 8.060 144.710 8.280 ;
        RECT 147.460 8.210 147.870 8.640 ;
        RECT 148.260 8.540 148.710 8.640 ;
        RECT 149.920 8.880 150.370 8.990 ;
        RECT 151.770 8.880 152.220 8.990 ;
        RECT 149.920 8.640 152.220 8.880 ;
        RECT 149.920 8.540 150.370 8.640 ;
        RECT 150.760 8.210 151.170 8.640 ;
        RECT 151.770 8.570 152.220 8.640 ;
        RECT 153.170 8.880 153.620 8.960 ;
        RECT 154.220 8.880 154.630 9.320 ;
        RECT 155.020 8.880 155.470 8.990 ;
        RECT 153.170 8.640 155.470 8.880 ;
        RECT 153.170 8.540 153.620 8.640 ;
        RECT 155.020 8.540 155.470 8.640 ;
        RECT 156.660 8.880 157.110 8.990 ;
        RECT 157.500 8.880 157.910 9.320 ;
        RECT 160.680 9.050 161.130 9.330 ;
        RECT 164.500 9.050 164.950 9.330 ;
        RECT 174.180 9.330 175.710 9.540 ;
        RECT 176.090 9.450 176.540 9.540 ;
        RECT 176.920 9.330 178.450 9.540 ;
        RECT 158.510 8.880 158.960 8.960 ;
        RECT 156.660 8.640 158.960 8.880 ;
        RECT 156.660 8.540 157.110 8.640 ;
        RECT 158.510 8.540 158.960 8.640 ;
        RECT 159.910 8.880 160.360 8.990 ;
        RECT 161.760 8.880 162.210 8.990 ;
        RECT 159.910 8.640 162.210 8.880 ;
        RECT 159.910 8.570 160.360 8.640 ;
        RECT 143.160 8.010 143.610 8.060 ;
        RECT 141.520 7.720 143.610 8.010 ;
        RECT 141.520 7.670 141.970 7.720 ;
        RECT 124.770 7.090 125.220 7.160 ;
        RECT 122.920 6.850 125.220 7.090 ;
        RECT 122.920 6.740 123.370 6.850 ;
        RECT 124.770 6.740 125.220 6.850 ;
        RECT 126.170 7.090 126.620 7.190 ;
        RECT 128.020 7.090 128.470 7.190 ;
        RECT 126.170 6.850 128.470 7.090 ;
        RECT 126.170 6.770 126.620 6.850 ;
        RECT 106.680 6.190 108.210 6.400 ;
        RECT 108.590 6.190 109.040 6.280 ;
        RECT 109.420 6.190 110.950 6.400 ;
        RECT 120.180 6.400 120.630 6.680 ;
        RECT 124.000 6.400 124.450 6.680 ;
        RECT 127.220 6.410 127.630 6.850 ;
        RECT 128.020 6.740 128.470 6.850 ;
        RECT 129.660 7.090 130.110 7.190 ;
        RECT 131.510 7.090 131.960 7.190 ;
        RECT 129.660 6.850 131.960 7.090 ;
        RECT 129.660 6.740 130.110 6.850 ;
        RECT 130.500 6.410 130.910 6.850 ;
        RECT 131.510 6.770 131.960 6.850 ;
        RECT 132.910 7.090 133.360 7.160 ;
        RECT 133.960 7.090 134.370 7.520 ;
        RECT 134.760 7.090 135.210 7.190 ;
        RECT 132.910 6.850 135.210 7.090 ;
        RECT 132.910 6.740 133.360 6.850 ;
        RECT 134.760 6.740 135.210 6.850 ;
        RECT 136.420 7.090 136.870 7.190 ;
        RECT 137.260 7.090 137.670 7.520 ;
        RECT 140.420 7.450 141.970 7.670 ;
        RECT 142.350 7.660 142.780 7.720 ;
        RECT 143.160 7.670 143.610 7.720 ;
        RECT 144.210 7.670 144.710 8.060 ;
        RECT 143.160 7.450 144.710 7.670 ;
        RECT 153.920 8.060 155.470 8.280 ;
        RECT 153.920 7.670 154.420 8.060 ;
        RECT 155.020 8.010 155.470 8.060 ;
        RECT 155.850 8.010 156.280 8.070 ;
        RECT 156.660 8.060 158.210 8.280 ;
        RECT 160.960 8.210 161.370 8.640 ;
        RECT 161.760 8.540 162.210 8.640 ;
        RECT 163.420 8.880 163.870 8.990 ;
        RECT 165.270 8.880 165.720 8.990 ;
        RECT 163.420 8.640 165.720 8.880 ;
        RECT 163.420 8.540 163.870 8.640 ;
        RECT 164.260 8.210 164.670 8.640 ;
        RECT 165.270 8.570 165.720 8.640 ;
        RECT 166.670 8.880 167.120 8.960 ;
        RECT 167.720 8.880 168.130 9.320 ;
        RECT 168.520 8.880 168.970 8.990 ;
        RECT 166.670 8.640 168.970 8.880 ;
        RECT 166.670 8.540 167.120 8.640 ;
        RECT 168.520 8.540 168.970 8.640 ;
        RECT 170.160 8.880 170.610 8.990 ;
        RECT 171.000 8.880 171.410 9.320 ;
        RECT 174.180 9.050 174.630 9.330 ;
        RECT 178.000 9.050 178.450 9.330 ;
        RECT 187.680 9.330 189.210 9.540 ;
        RECT 189.590 9.450 190.040 9.540 ;
        RECT 190.420 9.330 191.950 9.540 ;
        RECT 172.010 8.880 172.460 8.960 ;
        RECT 170.160 8.640 172.460 8.880 ;
        RECT 170.160 8.540 170.610 8.640 ;
        RECT 172.010 8.540 172.460 8.640 ;
        RECT 173.410 8.880 173.860 8.990 ;
        RECT 175.260 8.880 175.710 8.990 ;
        RECT 173.410 8.640 175.710 8.880 ;
        RECT 173.410 8.570 173.860 8.640 ;
        RECT 156.660 8.010 157.110 8.060 ;
        RECT 155.020 7.720 157.110 8.010 ;
        RECT 155.020 7.670 155.470 7.720 ;
        RECT 138.270 7.090 138.720 7.160 ;
        RECT 136.420 6.850 138.720 7.090 ;
        RECT 136.420 6.740 136.870 6.850 ;
        RECT 138.270 6.740 138.720 6.850 ;
        RECT 139.670 7.090 140.120 7.190 ;
        RECT 141.520 7.090 141.970 7.190 ;
        RECT 139.670 6.850 141.970 7.090 ;
        RECT 139.670 6.770 140.120 6.850 ;
        RECT 120.180 6.190 121.710 6.400 ;
        RECT 122.090 6.190 122.540 6.280 ;
        RECT 122.920 6.190 124.450 6.400 ;
        RECT 133.680 6.400 134.130 6.680 ;
        RECT 137.500 6.400 137.950 6.680 ;
        RECT 140.720 6.410 141.130 6.850 ;
        RECT 141.520 6.740 141.970 6.850 ;
        RECT 143.160 7.090 143.610 7.190 ;
        RECT 145.010 7.090 145.460 7.190 ;
        RECT 143.160 6.850 145.460 7.090 ;
        RECT 143.160 6.740 143.610 6.850 ;
        RECT 144.000 6.410 144.410 6.850 ;
        RECT 145.010 6.770 145.460 6.850 ;
        RECT 146.410 7.090 146.860 7.160 ;
        RECT 147.460 7.090 147.870 7.520 ;
        RECT 148.260 7.090 148.710 7.190 ;
        RECT 146.410 6.850 148.710 7.090 ;
        RECT 146.410 6.740 146.860 6.850 ;
        RECT 148.260 6.740 148.710 6.850 ;
        RECT 149.920 7.090 150.370 7.190 ;
        RECT 150.760 7.090 151.170 7.520 ;
        RECT 153.920 7.450 155.470 7.670 ;
        RECT 155.850 7.660 156.280 7.720 ;
        RECT 156.660 7.670 157.110 7.720 ;
        RECT 157.710 7.670 158.210 8.060 ;
        RECT 156.660 7.450 158.210 7.670 ;
        RECT 167.420 8.060 168.970 8.280 ;
        RECT 167.420 7.670 167.920 8.060 ;
        RECT 168.520 8.010 168.970 8.060 ;
        RECT 169.350 8.010 169.780 8.070 ;
        RECT 170.160 8.060 171.710 8.280 ;
        RECT 174.460 8.210 174.870 8.640 ;
        RECT 175.260 8.540 175.710 8.640 ;
        RECT 176.920 8.880 177.370 8.990 ;
        RECT 178.770 8.880 179.220 8.990 ;
        RECT 176.920 8.640 179.220 8.880 ;
        RECT 176.920 8.540 177.370 8.640 ;
        RECT 177.760 8.210 178.170 8.640 ;
        RECT 178.770 8.570 179.220 8.640 ;
        RECT 180.170 8.880 180.620 8.960 ;
        RECT 181.220 8.880 181.630 9.320 ;
        RECT 182.020 8.880 182.470 8.990 ;
        RECT 180.170 8.640 182.470 8.880 ;
        RECT 180.170 8.540 180.620 8.640 ;
        RECT 182.020 8.540 182.470 8.640 ;
        RECT 183.660 8.880 184.110 8.990 ;
        RECT 184.500 8.880 184.910 9.320 ;
        RECT 187.680 9.050 188.130 9.330 ;
        RECT 191.500 9.050 191.950 9.330 ;
        RECT 201.180 9.330 202.710 9.540 ;
        RECT 203.090 9.450 203.540 9.540 ;
        RECT 203.920 9.330 205.450 9.540 ;
        RECT 185.510 8.880 185.960 8.960 ;
        RECT 183.660 8.640 185.960 8.880 ;
        RECT 183.660 8.540 184.110 8.640 ;
        RECT 185.510 8.540 185.960 8.640 ;
        RECT 186.910 8.880 187.360 8.990 ;
        RECT 188.760 8.880 189.210 8.990 ;
        RECT 186.910 8.640 189.210 8.880 ;
        RECT 186.910 8.570 187.360 8.640 ;
        RECT 170.160 8.010 170.610 8.060 ;
        RECT 168.520 7.720 170.610 8.010 ;
        RECT 168.520 7.670 168.970 7.720 ;
        RECT 151.770 7.090 152.220 7.160 ;
        RECT 149.920 6.850 152.220 7.090 ;
        RECT 149.920 6.740 150.370 6.850 ;
        RECT 151.770 6.740 152.220 6.850 ;
        RECT 153.170 7.090 153.620 7.190 ;
        RECT 155.020 7.090 155.470 7.190 ;
        RECT 153.170 6.850 155.470 7.090 ;
        RECT 153.170 6.770 153.620 6.850 ;
        RECT 133.680 6.190 135.210 6.400 ;
        RECT 135.590 6.190 136.040 6.280 ;
        RECT 136.420 6.190 137.950 6.400 ;
        RECT 147.180 6.400 147.630 6.680 ;
        RECT 151.000 6.400 151.450 6.680 ;
        RECT 154.220 6.410 154.630 6.850 ;
        RECT 155.020 6.740 155.470 6.850 ;
        RECT 156.660 7.090 157.110 7.190 ;
        RECT 158.510 7.090 158.960 7.190 ;
        RECT 156.660 6.850 158.960 7.090 ;
        RECT 156.660 6.740 157.110 6.850 ;
        RECT 157.500 6.410 157.910 6.850 ;
        RECT 158.510 6.770 158.960 6.850 ;
        RECT 159.910 7.090 160.360 7.160 ;
        RECT 160.960 7.090 161.370 7.520 ;
        RECT 161.760 7.090 162.210 7.190 ;
        RECT 159.910 6.850 162.210 7.090 ;
        RECT 159.910 6.740 160.360 6.850 ;
        RECT 161.760 6.740 162.210 6.850 ;
        RECT 163.420 7.090 163.870 7.190 ;
        RECT 164.260 7.090 164.670 7.520 ;
        RECT 167.420 7.450 168.970 7.670 ;
        RECT 169.350 7.660 169.780 7.720 ;
        RECT 170.160 7.670 170.610 7.720 ;
        RECT 171.210 7.670 171.710 8.060 ;
        RECT 170.160 7.450 171.710 7.670 ;
        RECT 180.920 8.060 182.470 8.280 ;
        RECT 180.920 7.670 181.420 8.060 ;
        RECT 182.020 8.010 182.470 8.060 ;
        RECT 182.850 8.010 183.280 8.070 ;
        RECT 183.660 8.060 185.210 8.280 ;
        RECT 187.960 8.210 188.370 8.640 ;
        RECT 188.760 8.540 189.210 8.640 ;
        RECT 190.420 8.880 190.870 8.990 ;
        RECT 192.270 8.880 192.720 8.990 ;
        RECT 190.420 8.640 192.720 8.880 ;
        RECT 190.420 8.540 190.870 8.640 ;
        RECT 191.260 8.210 191.670 8.640 ;
        RECT 192.270 8.570 192.720 8.640 ;
        RECT 193.670 8.880 194.120 8.960 ;
        RECT 194.720 8.880 195.130 9.320 ;
        RECT 195.520 8.880 195.970 8.990 ;
        RECT 193.670 8.640 195.970 8.880 ;
        RECT 193.670 8.540 194.120 8.640 ;
        RECT 195.520 8.540 195.970 8.640 ;
        RECT 197.160 8.880 197.610 8.990 ;
        RECT 198.000 8.880 198.410 9.320 ;
        RECT 201.180 9.050 201.630 9.330 ;
        RECT 205.000 9.050 205.450 9.330 ;
        RECT 214.680 9.330 216.210 9.540 ;
        RECT 216.590 9.450 217.030 9.540 ;
        RECT 199.010 8.880 199.460 8.960 ;
        RECT 197.160 8.640 199.460 8.880 ;
        RECT 197.160 8.540 197.610 8.640 ;
        RECT 199.010 8.540 199.460 8.640 ;
        RECT 200.410 8.880 200.860 8.990 ;
        RECT 202.260 8.880 202.710 8.990 ;
        RECT 200.410 8.640 202.710 8.880 ;
        RECT 200.410 8.570 200.860 8.640 ;
        RECT 183.660 8.010 184.110 8.060 ;
        RECT 182.020 7.720 184.110 8.010 ;
        RECT 182.020 7.670 182.470 7.720 ;
        RECT 165.270 7.090 165.720 7.160 ;
        RECT 163.420 6.850 165.720 7.090 ;
        RECT 163.420 6.740 163.870 6.850 ;
        RECT 165.270 6.740 165.720 6.850 ;
        RECT 166.670 7.090 167.120 7.190 ;
        RECT 168.520 7.090 168.970 7.190 ;
        RECT 166.670 6.850 168.970 7.090 ;
        RECT 166.670 6.770 167.120 6.850 ;
        RECT 147.180 6.190 148.710 6.400 ;
        RECT 149.090 6.190 149.540 6.280 ;
        RECT 149.920 6.190 151.450 6.400 ;
        RECT 160.680 6.400 161.130 6.680 ;
        RECT 164.500 6.400 164.950 6.680 ;
        RECT 167.720 6.410 168.130 6.850 ;
        RECT 168.520 6.740 168.970 6.850 ;
        RECT 170.160 7.090 170.610 7.190 ;
        RECT 172.010 7.090 172.460 7.190 ;
        RECT 170.160 6.850 172.460 7.090 ;
        RECT 170.160 6.740 170.610 6.850 ;
        RECT 171.000 6.410 171.410 6.850 ;
        RECT 172.010 6.770 172.460 6.850 ;
        RECT 173.410 7.090 173.860 7.160 ;
        RECT 174.460 7.090 174.870 7.520 ;
        RECT 175.260 7.090 175.710 7.190 ;
        RECT 173.410 6.850 175.710 7.090 ;
        RECT 173.410 6.740 173.860 6.850 ;
        RECT 175.260 6.740 175.710 6.850 ;
        RECT 176.920 7.090 177.370 7.190 ;
        RECT 177.760 7.090 178.170 7.520 ;
        RECT 180.920 7.450 182.470 7.670 ;
        RECT 182.850 7.660 183.280 7.720 ;
        RECT 183.660 7.670 184.110 7.720 ;
        RECT 184.710 7.670 185.210 8.060 ;
        RECT 183.660 7.450 185.210 7.670 ;
        RECT 194.420 8.060 195.970 8.280 ;
        RECT 194.420 7.670 194.920 8.060 ;
        RECT 195.520 8.010 195.970 8.060 ;
        RECT 196.350 8.010 196.780 8.070 ;
        RECT 197.160 8.060 198.710 8.280 ;
        RECT 201.460 8.210 201.870 8.640 ;
        RECT 202.260 8.540 202.710 8.640 ;
        RECT 203.920 8.880 204.370 8.990 ;
        RECT 205.770 8.880 206.220 8.990 ;
        RECT 203.920 8.640 206.220 8.880 ;
        RECT 203.920 8.540 204.370 8.640 ;
        RECT 204.760 8.210 205.170 8.640 ;
        RECT 205.770 8.570 206.220 8.640 ;
        RECT 207.170 8.880 207.620 8.960 ;
        RECT 208.220 8.880 208.630 9.320 ;
        RECT 209.020 8.880 209.470 8.990 ;
        RECT 207.170 8.640 209.470 8.880 ;
        RECT 207.170 8.540 207.620 8.640 ;
        RECT 209.020 8.540 209.470 8.640 ;
        RECT 210.660 8.880 211.110 8.990 ;
        RECT 211.500 8.880 211.910 9.320 ;
        RECT 214.680 9.050 215.130 9.330 ;
        RECT 212.510 8.880 212.960 8.960 ;
        RECT 210.660 8.640 212.960 8.880 ;
        RECT 210.660 8.540 211.110 8.640 ;
        RECT 212.510 8.540 212.960 8.640 ;
        RECT 213.910 8.880 214.360 8.990 ;
        RECT 215.760 8.880 216.210 8.990 ;
        RECT 213.910 8.640 216.210 8.880 ;
        RECT 213.910 8.570 214.360 8.640 ;
        RECT 197.160 8.010 197.610 8.060 ;
        RECT 195.520 7.720 197.610 8.010 ;
        RECT 195.520 7.670 195.970 7.720 ;
        RECT 178.770 7.090 179.220 7.160 ;
        RECT 176.920 6.850 179.220 7.090 ;
        RECT 176.920 6.740 177.370 6.850 ;
        RECT 178.770 6.740 179.220 6.850 ;
        RECT 180.170 7.090 180.620 7.190 ;
        RECT 182.020 7.090 182.470 7.190 ;
        RECT 180.170 6.850 182.470 7.090 ;
        RECT 180.170 6.770 180.620 6.850 ;
        RECT 160.680 6.190 162.210 6.400 ;
        RECT 162.590 6.190 163.040 6.280 ;
        RECT 163.420 6.190 164.950 6.400 ;
        RECT 174.180 6.400 174.630 6.680 ;
        RECT 178.000 6.400 178.450 6.680 ;
        RECT 181.220 6.410 181.630 6.850 ;
        RECT 182.020 6.740 182.470 6.850 ;
        RECT 183.660 7.090 184.110 7.190 ;
        RECT 185.510 7.090 185.960 7.190 ;
        RECT 183.660 6.850 185.960 7.090 ;
        RECT 183.660 6.740 184.110 6.850 ;
        RECT 184.500 6.410 184.910 6.850 ;
        RECT 185.510 6.770 185.960 6.850 ;
        RECT 186.910 7.090 187.360 7.160 ;
        RECT 187.960 7.090 188.370 7.520 ;
        RECT 188.760 7.090 189.210 7.190 ;
        RECT 186.910 6.850 189.210 7.090 ;
        RECT 186.910 6.740 187.360 6.850 ;
        RECT 188.760 6.740 189.210 6.850 ;
        RECT 190.420 7.090 190.870 7.190 ;
        RECT 191.260 7.090 191.670 7.520 ;
        RECT 194.420 7.450 195.970 7.670 ;
        RECT 196.350 7.660 196.780 7.720 ;
        RECT 197.160 7.670 197.610 7.720 ;
        RECT 198.210 7.670 198.710 8.060 ;
        RECT 197.160 7.450 198.710 7.670 ;
        RECT 207.920 8.060 209.470 8.280 ;
        RECT 207.920 7.670 208.420 8.060 ;
        RECT 209.020 8.010 209.470 8.060 ;
        RECT 209.850 8.010 210.280 8.070 ;
        RECT 210.660 8.060 212.210 8.280 ;
        RECT 214.960 8.210 215.370 8.640 ;
        RECT 215.760 8.540 216.210 8.640 ;
        RECT 210.660 8.010 211.110 8.060 ;
        RECT 209.020 7.720 211.110 8.010 ;
        RECT 209.020 7.670 209.470 7.720 ;
        RECT 192.270 7.090 192.720 7.160 ;
        RECT 190.420 6.850 192.720 7.090 ;
        RECT 190.420 6.740 190.870 6.850 ;
        RECT 192.270 6.740 192.720 6.850 ;
        RECT 193.670 7.090 194.120 7.190 ;
        RECT 195.520 7.090 195.970 7.190 ;
        RECT 193.670 6.850 195.970 7.090 ;
        RECT 193.670 6.770 194.120 6.850 ;
        RECT 174.180 6.190 175.710 6.400 ;
        RECT 176.090 6.190 176.540 6.280 ;
        RECT 176.920 6.190 178.450 6.400 ;
        RECT 187.680 6.400 188.130 6.680 ;
        RECT 191.500 6.400 191.950 6.680 ;
        RECT 194.720 6.410 195.130 6.850 ;
        RECT 195.520 6.740 195.970 6.850 ;
        RECT 197.160 7.090 197.610 7.190 ;
        RECT 199.010 7.090 199.460 7.190 ;
        RECT 197.160 6.850 199.460 7.090 ;
        RECT 197.160 6.740 197.610 6.850 ;
        RECT 198.000 6.410 198.410 6.850 ;
        RECT 199.010 6.770 199.460 6.850 ;
        RECT 200.410 7.090 200.860 7.160 ;
        RECT 201.460 7.090 201.870 7.520 ;
        RECT 202.260 7.090 202.710 7.190 ;
        RECT 200.410 6.850 202.710 7.090 ;
        RECT 200.410 6.740 200.860 6.850 ;
        RECT 202.260 6.740 202.710 6.850 ;
        RECT 203.920 7.090 204.370 7.190 ;
        RECT 204.760 7.090 205.170 7.520 ;
        RECT 207.920 7.450 209.470 7.670 ;
        RECT 209.850 7.660 210.280 7.720 ;
        RECT 210.660 7.670 211.110 7.720 ;
        RECT 211.710 7.670 212.210 8.060 ;
        RECT 210.660 7.450 212.210 7.670 ;
        RECT 205.770 7.090 206.220 7.160 ;
        RECT 203.920 6.850 206.220 7.090 ;
        RECT 203.920 6.740 204.370 6.850 ;
        RECT 205.770 6.740 206.220 6.850 ;
        RECT 207.170 7.090 207.620 7.190 ;
        RECT 209.020 7.090 209.470 7.190 ;
        RECT 207.170 6.850 209.470 7.090 ;
        RECT 207.170 6.770 207.620 6.850 ;
        RECT 187.680 6.190 189.210 6.400 ;
        RECT 189.590 6.190 190.040 6.280 ;
        RECT 190.420 6.190 191.950 6.400 ;
        RECT 201.180 6.400 201.630 6.680 ;
        RECT 205.000 6.400 205.450 6.680 ;
        RECT 208.220 6.410 208.630 6.850 ;
        RECT 209.020 6.740 209.470 6.850 ;
        RECT 210.660 7.090 211.110 7.190 ;
        RECT 212.510 7.090 212.960 7.190 ;
        RECT 210.660 6.850 212.960 7.090 ;
        RECT 210.660 6.740 211.110 6.850 ;
        RECT 211.500 6.410 211.910 6.850 ;
        RECT 212.510 6.770 212.960 6.850 ;
        RECT 213.910 7.090 214.360 7.160 ;
        RECT 214.960 7.090 215.370 7.520 ;
        RECT 215.760 7.090 216.210 7.190 ;
        RECT 213.910 6.850 216.210 7.090 ;
        RECT 213.910 6.740 214.360 6.850 ;
        RECT 215.760 6.740 216.210 6.850 ;
        RECT 201.180 6.190 202.710 6.400 ;
        RECT 203.090 6.190 203.540 6.280 ;
        RECT 203.920 6.190 205.450 6.400 ;
        RECT 214.680 6.400 215.130 6.680 ;
        RECT 214.680 6.190 216.210 6.400 ;
        RECT 216.590 6.190 217.030 6.280 ;
        RECT 13.260 5.930 15.370 6.190 ;
        RECT 26.760 5.930 28.870 6.190 ;
        RECT 40.260 5.930 42.370 6.190 ;
        RECT 53.760 5.930 55.870 6.190 ;
        RECT 67.260 5.930 69.370 6.190 ;
        RECT 80.760 5.930 82.870 6.190 ;
        RECT 94.260 5.930 96.370 6.190 ;
        RECT 107.760 5.930 109.870 6.190 ;
        RECT 121.260 5.930 123.370 6.190 ;
        RECT 134.760 5.930 136.870 6.190 ;
        RECT 148.260 5.930 150.370 6.190 ;
        RECT 161.760 5.930 163.870 6.190 ;
        RECT 175.260 5.930 177.370 6.190 ;
        RECT 188.760 5.930 190.870 6.190 ;
        RECT 202.260 5.930 204.370 6.190 ;
        RECT 215.760 6.130 217.030 6.190 ;
        RECT 215.760 5.940 217.240 6.130 ;
        RECT 215.760 5.930 217.030 5.940 ;
        RECT 12.180 5.720 13.710 5.930 ;
        RECT 14.090 5.840 14.540 5.930 ;
        RECT 14.920 5.720 16.450 5.930 ;
        RECT 1.420 5.270 1.870 5.380 ;
        RECT 3.270 5.270 3.720 5.380 ;
        RECT 1.420 5.030 3.720 5.270 ;
        RECT 1.420 4.930 1.870 5.030 ;
        RECT 2.260 4.600 2.670 5.030 ;
        RECT 3.270 4.960 3.720 5.030 ;
        RECT 4.670 5.270 5.120 5.350 ;
        RECT 5.720 5.270 6.130 5.710 ;
        RECT 6.520 5.270 6.970 5.380 ;
        RECT 4.670 5.030 6.970 5.270 ;
        RECT 4.670 4.930 5.120 5.030 ;
        RECT 6.520 4.930 6.970 5.030 ;
        RECT 8.160 5.270 8.610 5.380 ;
        RECT 9.000 5.270 9.410 5.710 ;
        RECT 12.180 5.440 12.630 5.720 ;
        RECT 16.000 5.440 16.450 5.720 ;
        RECT 25.680 5.720 27.210 5.930 ;
        RECT 27.590 5.840 28.040 5.930 ;
        RECT 28.420 5.720 29.950 5.930 ;
        RECT 10.010 5.270 10.460 5.350 ;
        RECT 8.160 5.030 10.460 5.270 ;
        RECT 8.160 4.930 8.610 5.030 ;
        RECT 10.010 4.930 10.460 5.030 ;
        RECT 11.410 5.270 11.860 5.380 ;
        RECT 13.260 5.270 13.710 5.380 ;
        RECT 11.410 5.030 13.710 5.270 ;
        RECT 11.410 4.960 11.860 5.030 ;
        RECT 5.420 4.450 6.970 4.670 ;
        RECT 5.420 4.060 5.920 4.450 ;
        RECT 6.520 4.400 6.970 4.450 ;
        RECT 7.350 4.400 7.780 4.460 ;
        RECT 8.160 4.450 9.710 4.670 ;
        RECT 12.460 4.600 12.870 5.030 ;
        RECT 13.260 4.930 13.710 5.030 ;
        RECT 14.920 5.270 15.370 5.380 ;
        RECT 16.770 5.270 17.220 5.380 ;
        RECT 14.920 5.030 17.220 5.270 ;
        RECT 14.920 4.930 15.370 5.030 ;
        RECT 15.760 4.600 16.170 5.030 ;
        RECT 16.770 4.960 17.220 5.030 ;
        RECT 18.170 5.270 18.620 5.350 ;
        RECT 19.220 5.270 19.630 5.710 ;
        RECT 20.020 5.270 20.470 5.380 ;
        RECT 18.170 5.030 20.470 5.270 ;
        RECT 18.170 4.930 18.620 5.030 ;
        RECT 20.020 4.930 20.470 5.030 ;
        RECT 21.660 5.270 22.110 5.380 ;
        RECT 22.500 5.270 22.910 5.710 ;
        RECT 25.680 5.440 26.130 5.720 ;
        RECT 29.500 5.440 29.950 5.720 ;
        RECT 39.180 5.720 40.710 5.930 ;
        RECT 41.090 5.840 41.540 5.930 ;
        RECT 41.920 5.720 43.450 5.930 ;
        RECT 23.510 5.270 23.960 5.350 ;
        RECT 21.660 5.030 23.960 5.270 ;
        RECT 21.660 4.930 22.110 5.030 ;
        RECT 23.510 4.930 23.960 5.030 ;
        RECT 24.910 5.270 25.360 5.380 ;
        RECT 26.760 5.270 27.210 5.380 ;
        RECT 24.910 5.030 27.210 5.270 ;
        RECT 24.910 4.960 25.360 5.030 ;
        RECT 8.160 4.400 8.610 4.450 ;
        RECT 6.520 4.110 8.610 4.400 ;
        RECT 6.520 4.060 6.970 4.110 ;
        RECT 1.420 3.480 1.870 3.580 ;
        RECT 2.260 3.480 2.670 3.910 ;
        RECT 5.420 3.840 6.970 4.060 ;
        RECT 7.350 4.050 7.780 4.110 ;
        RECT 8.160 4.060 8.610 4.110 ;
        RECT 9.210 4.060 9.710 4.450 ;
        RECT 8.160 3.840 9.710 4.060 ;
        RECT 18.920 4.450 20.470 4.670 ;
        RECT 18.920 4.060 19.420 4.450 ;
        RECT 20.020 4.400 20.470 4.450 ;
        RECT 20.850 4.400 21.280 4.460 ;
        RECT 21.660 4.450 23.210 4.670 ;
        RECT 25.960 4.600 26.370 5.030 ;
        RECT 26.760 4.930 27.210 5.030 ;
        RECT 28.420 5.270 28.870 5.380 ;
        RECT 30.270 5.270 30.720 5.380 ;
        RECT 28.420 5.030 30.720 5.270 ;
        RECT 28.420 4.930 28.870 5.030 ;
        RECT 29.260 4.600 29.670 5.030 ;
        RECT 30.270 4.960 30.720 5.030 ;
        RECT 31.670 5.270 32.120 5.350 ;
        RECT 32.720 5.270 33.130 5.710 ;
        RECT 33.520 5.270 33.970 5.380 ;
        RECT 31.670 5.030 33.970 5.270 ;
        RECT 31.670 4.930 32.120 5.030 ;
        RECT 33.520 4.930 33.970 5.030 ;
        RECT 35.160 5.270 35.610 5.380 ;
        RECT 36.000 5.270 36.410 5.710 ;
        RECT 39.180 5.440 39.630 5.720 ;
        RECT 43.000 5.440 43.450 5.720 ;
        RECT 52.680 5.720 54.210 5.930 ;
        RECT 54.590 5.840 55.040 5.930 ;
        RECT 55.420 5.720 56.950 5.930 ;
        RECT 37.010 5.270 37.460 5.350 ;
        RECT 35.160 5.030 37.460 5.270 ;
        RECT 35.160 4.930 35.610 5.030 ;
        RECT 37.010 4.930 37.460 5.030 ;
        RECT 38.410 5.270 38.860 5.380 ;
        RECT 40.260 5.270 40.710 5.380 ;
        RECT 38.410 5.030 40.710 5.270 ;
        RECT 38.410 4.960 38.860 5.030 ;
        RECT 21.660 4.400 22.110 4.450 ;
        RECT 20.020 4.110 22.110 4.400 ;
        RECT 20.020 4.060 20.470 4.110 ;
        RECT 3.270 3.480 3.720 3.550 ;
        RECT 1.420 3.240 3.720 3.480 ;
        RECT 1.420 3.130 1.870 3.240 ;
        RECT 3.270 3.130 3.720 3.240 ;
        RECT 4.670 3.480 5.120 3.580 ;
        RECT 6.520 3.480 6.970 3.580 ;
        RECT 4.670 3.240 6.970 3.480 ;
        RECT 4.670 3.160 5.120 3.240 ;
        RECT 5.720 2.800 6.130 3.240 ;
        RECT 6.520 3.130 6.970 3.240 ;
        RECT 8.160 3.480 8.610 3.580 ;
        RECT 10.010 3.480 10.460 3.580 ;
        RECT 8.160 3.240 10.460 3.480 ;
        RECT 8.160 3.130 8.610 3.240 ;
        RECT 9.000 2.800 9.410 3.240 ;
        RECT 10.010 3.160 10.460 3.240 ;
        RECT 11.410 3.480 11.860 3.550 ;
        RECT 12.460 3.480 12.870 3.910 ;
        RECT 13.260 3.480 13.710 3.580 ;
        RECT 11.410 3.240 13.710 3.480 ;
        RECT 11.410 3.130 11.860 3.240 ;
        RECT 13.260 3.130 13.710 3.240 ;
        RECT 14.920 3.480 15.370 3.580 ;
        RECT 15.760 3.480 16.170 3.910 ;
        RECT 18.920 3.840 20.470 4.060 ;
        RECT 20.850 4.050 21.280 4.110 ;
        RECT 21.660 4.060 22.110 4.110 ;
        RECT 22.710 4.060 23.210 4.450 ;
        RECT 21.660 3.840 23.210 4.060 ;
        RECT 32.420 4.450 33.970 4.670 ;
        RECT 32.420 4.060 32.920 4.450 ;
        RECT 33.520 4.400 33.970 4.450 ;
        RECT 34.350 4.400 34.780 4.460 ;
        RECT 35.160 4.450 36.710 4.670 ;
        RECT 39.460 4.600 39.870 5.030 ;
        RECT 40.260 4.930 40.710 5.030 ;
        RECT 41.920 5.270 42.370 5.380 ;
        RECT 43.770 5.270 44.220 5.380 ;
        RECT 41.920 5.030 44.220 5.270 ;
        RECT 41.920 4.930 42.370 5.030 ;
        RECT 42.760 4.600 43.170 5.030 ;
        RECT 43.770 4.960 44.220 5.030 ;
        RECT 45.170 5.270 45.620 5.350 ;
        RECT 46.220 5.270 46.630 5.710 ;
        RECT 47.020 5.270 47.470 5.380 ;
        RECT 45.170 5.030 47.470 5.270 ;
        RECT 45.170 4.930 45.620 5.030 ;
        RECT 47.020 4.930 47.470 5.030 ;
        RECT 48.660 5.270 49.110 5.380 ;
        RECT 49.500 5.270 49.910 5.710 ;
        RECT 52.680 5.440 53.130 5.720 ;
        RECT 56.500 5.440 56.950 5.720 ;
        RECT 66.180 5.720 67.710 5.930 ;
        RECT 68.090 5.840 68.540 5.930 ;
        RECT 68.920 5.720 70.450 5.930 ;
        RECT 50.510 5.270 50.960 5.350 ;
        RECT 48.660 5.030 50.960 5.270 ;
        RECT 48.660 4.930 49.110 5.030 ;
        RECT 50.510 4.930 50.960 5.030 ;
        RECT 51.910 5.270 52.360 5.380 ;
        RECT 53.760 5.270 54.210 5.380 ;
        RECT 51.910 5.030 54.210 5.270 ;
        RECT 51.910 4.960 52.360 5.030 ;
        RECT 35.160 4.400 35.610 4.450 ;
        RECT 33.520 4.110 35.610 4.400 ;
        RECT 33.520 4.060 33.970 4.110 ;
        RECT 16.770 3.480 17.220 3.550 ;
        RECT 14.920 3.240 17.220 3.480 ;
        RECT 14.920 3.130 15.370 3.240 ;
        RECT 16.770 3.130 17.220 3.240 ;
        RECT 18.170 3.480 18.620 3.580 ;
        RECT 20.020 3.480 20.470 3.580 ;
        RECT 18.170 3.240 20.470 3.480 ;
        RECT 18.170 3.160 18.620 3.240 ;
        RECT 12.180 2.790 12.630 3.070 ;
        RECT 16.000 2.790 16.450 3.070 ;
        RECT 19.220 2.800 19.630 3.240 ;
        RECT 20.020 3.130 20.470 3.240 ;
        RECT 21.660 3.480 22.110 3.580 ;
        RECT 23.510 3.480 23.960 3.580 ;
        RECT 21.660 3.240 23.960 3.480 ;
        RECT 21.660 3.130 22.110 3.240 ;
        RECT 22.500 2.800 22.910 3.240 ;
        RECT 23.510 3.160 23.960 3.240 ;
        RECT 24.910 3.480 25.360 3.550 ;
        RECT 25.960 3.480 26.370 3.910 ;
        RECT 26.760 3.480 27.210 3.580 ;
        RECT 24.910 3.240 27.210 3.480 ;
        RECT 24.910 3.130 25.360 3.240 ;
        RECT 26.760 3.130 27.210 3.240 ;
        RECT 28.420 3.480 28.870 3.580 ;
        RECT 29.260 3.480 29.670 3.910 ;
        RECT 32.420 3.840 33.970 4.060 ;
        RECT 34.350 4.050 34.780 4.110 ;
        RECT 35.160 4.060 35.610 4.110 ;
        RECT 36.210 4.060 36.710 4.450 ;
        RECT 35.160 3.840 36.710 4.060 ;
        RECT 45.920 4.450 47.470 4.670 ;
        RECT 45.920 4.060 46.420 4.450 ;
        RECT 47.020 4.400 47.470 4.450 ;
        RECT 47.850 4.400 48.280 4.460 ;
        RECT 48.660 4.450 50.210 4.670 ;
        RECT 52.960 4.600 53.370 5.030 ;
        RECT 53.760 4.930 54.210 5.030 ;
        RECT 55.420 5.270 55.870 5.380 ;
        RECT 57.270 5.270 57.720 5.380 ;
        RECT 55.420 5.030 57.720 5.270 ;
        RECT 55.420 4.930 55.870 5.030 ;
        RECT 56.260 4.600 56.670 5.030 ;
        RECT 57.270 4.960 57.720 5.030 ;
        RECT 58.670 5.270 59.120 5.350 ;
        RECT 59.720 5.270 60.130 5.710 ;
        RECT 60.520 5.270 60.970 5.380 ;
        RECT 58.670 5.030 60.970 5.270 ;
        RECT 58.670 4.930 59.120 5.030 ;
        RECT 60.520 4.930 60.970 5.030 ;
        RECT 62.160 5.270 62.610 5.380 ;
        RECT 63.000 5.270 63.410 5.710 ;
        RECT 66.180 5.440 66.630 5.720 ;
        RECT 70.000 5.440 70.450 5.720 ;
        RECT 79.680 5.720 81.210 5.930 ;
        RECT 81.590 5.840 82.040 5.930 ;
        RECT 82.420 5.720 83.950 5.930 ;
        RECT 64.010 5.270 64.460 5.350 ;
        RECT 62.160 5.030 64.460 5.270 ;
        RECT 62.160 4.930 62.610 5.030 ;
        RECT 64.010 4.930 64.460 5.030 ;
        RECT 65.410 5.270 65.860 5.380 ;
        RECT 67.260 5.270 67.710 5.380 ;
        RECT 65.410 5.030 67.710 5.270 ;
        RECT 65.410 4.960 65.860 5.030 ;
        RECT 48.660 4.400 49.110 4.450 ;
        RECT 47.020 4.110 49.110 4.400 ;
        RECT 47.020 4.060 47.470 4.110 ;
        RECT 30.270 3.480 30.720 3.550 ;
        RECT 28.420 3.240 30.720 3.480 ;
        RECT 28.420 3.130 28.870 3.240 ;
        RECT 30.270 3.130 30.720 3.240 ;
        RECT 31.670 3.480 32.120 3.580 ;
        RECT 33.520 3.480 33.970 3.580 ;
        RECT 31.670 3.240 33.970 3.480 ;
        RECT 31.670 3.160 32.120 3.240 ;
        RECT 12.180 2.580 13.710 2.790 ;
        RECT 14.090 2.580 14.540 2.670 ;
        RECT 14.920 2.580 16.450 2.790 ;
        RECT 25.680 2.790 26.130 3.070 ;
        RECT 29.500 2.790 29.950 3.070 ;
        RECT 32.720 2.800 33.130 3.240 ;
        RECT 33.520 3.130 33.970 3.240 ;
        RECT 35.160 3.480 35.610 3.580 ;
        RECT 37.010 3.480 37.460 3.580 ;
        RECT 35.160 3.240 37.460 3.480 ;
        RECT 35.160 3.130 35.610 3.240 ;
        RECT 36.000 2.800 36.410 3.240 ;
        RECT 37.010 3.160 37.460 3.240 ;
        RECT 38.410 3.480 38.860 3.550 ;
        RECT 39.460 3.480 39.870 3.910 ;
        RECT 40.260 3.480 40.710 3.580 ;
        RECT 38.410 3.240 40.710 3.480 ;
        RECT 38.410 3.130 38.860 3.240 ;
        RECT 40.260 3.130 40.710 3.240 ;
        RECT 41.920 3.480 42.370 3.580 ;
        RECT 42.760 3.480 43.170 3.910 ;
        RECT 45.920 3.840 47.470 4.060 ;
        RECT 47.850 4.050 48.280 4.110 ;
        RECT 48.660 4.060 49.110 4.110 ;
        RECT 49.710 4.060 50.210 4.450 ;
        RECT 48.660 3.840 50.210 4.060 ;
        RECT 59.420 4.450 60.970 4.670 ;
        RECT 59.420 4.060 59.920 4.450 ;
        RECT 60.520 4.400 60.970 4.450 ;
        RECT 61.350 4.400 61.780 4.460 ;
        RECT 62.160 4.450 63.710 4.670 ;
        RECT 66.460 4.600 66.870 5.030 ;
        RECT 67.260 4.930 67.710 5.030 ;
        RECT 68.920 5.270 69.370 5.380 ;
        RECT 70.770 5.270 71.220 5.380 ;
        RECT 68.920 5.030 71.220 5.270 ;
        RECT 68.920 4.930 69.370 5.030 ;
        RECT 69.760 4.600 70.170 5.030 ;
        RECT 70.770 4.960 71.220 5.030 ;
        RECT 72.170 5.270 72.620 5.350 ;
        RECT 73.220 5.270 73.630 5.710 ;
        RECT 74.020 5.270 74.470 5.380 ;
        RECT 72.170 5.030 74.470 5.270 ;
        RECT 72.170 4.930 72.620 5.030 ;
        RECT 74.020 4.930 74.470 5.030 ;
        RECT 75.660 5.270 76.110 5.380 ;
        RECT 76.500 5.270 76.910 5.710 ;
        RECT 79.680 5.440 80.130 5.720 ;
        RECT 83.500 5.440 83.950 5.720 ;
        RECT 93.180 5.720 94.710 5.930 ;
        RECT 95.090 5.840 95.540 5.930 ;
        RECT 95.920 5.720 97.450 5.930 ;
        RECT 77.510 5.270 77.960 5.350 ;
        RECT 75.660 5.030 77.960 5.270 ;
        RECT 75.660 4.930 76.110 5.030 ;
        RECT 77.510 4.930 77.960 5.030 ;
        RECT 78.910 5.270 79.360 5.380 ;
        RECT 80.760 5.270 81.210 5.380 ;
        RECT 78.910 5.030 81.210 5.270 ;
        RECT 78.910 4.960 79.360 5.030 ;
        RECT 62.160 4.400 62.610 4.450 ;
        RECT 60.520 4.110 62.610 4.400 ;
        RECT 60.520 4.060 60.970 4.110 ;
        RECT 43.770 3.480 44.220 3.550 ;
        RECT 41.920 3.240 44.220 3.480 ;
        RECT 41.920 3.130 42.370 3.240 ;
        RECT 43.770 3.130 44.220 3.240 ;
        RECT 45.170 3.480 45.620 3.580 ;
        RECT 47.020 3.480 47.470 3.580 ;
        RECT 45.170 3.240 47.470 3.480 ;
        RECT 45.170 3.160 45.620 3.240 ;
        RECT 25.680 2.580 27.210 2.790 ;
        RECT 27.590 2.580 28.040 2.670 ;
        RECT 28.420 2.580 29.950 2.790 ;
        RECT 39.180 2.790 39.630 3.070 ;
        RECT 43.000 2.790 43.450 3.070 ;
        RECT 46.220 2.800 46.630 3.240 ;
        RECT 47.020 3.130 47.470 3.240 ;
        RECT 48.660 3.480 49.110 3.580 ;
        RECT 50.510 3.480 50.960 3.580 ;
        RECT 48.660 3.240 50.960 3.480 ;
        RECT 48.660 3.130 49.110 3.240 ;
        RECT 49.500 2.800 49.910 3.240 ;
        RECT 50.510 3.160 50.960 3.240 ;
        RECT 51.910 3.480 52.360 3.550 ;
        RECT 52.960 3.480 53.370 3.910 ;
        RECT 53.760 3.480 54.210 3.580 ;
        RECT 51.910 3.240 54.210 3.480 ;
        RECT 51.910 3.130 52.360 3.240 ;
        RECT 53.760 3.130 54.210 3.240 ;
        RECT 55.420 3.480 55.870 3.580 ;
        RECT 56.260 3.480 56.670 3.910 ;
        RECT 59.420 3.840 60.970 4.060 ;
        RECT 61.350 4.050 61.780 4.110 ;
        RECT 62.160 4.060 62.610 4.110 ;
        RECT 63.210 4.060 63.710 4.450 ;
        RECT 62.160 3.840 63.710 4.060 ;
        RECT 72.920 4.450 74.470 4.670 ;
        RECT 72.920 4.060 73.420 4.450 ;
        RECT 74.020 4.400 74.470 4.450 ;
        RECT 74.850 4.400 75.280 4.460 ;
        RECT 75.660 4.450 77.210 4.670 ;
        RECT 79.960 4.600 80.370 5.030 ;
        RECT 80.760 4.930 81.210 5.030 ;
        RECT 82.420 5.270 82.870 5.380 ;
        RECT 84.270 5.270 84.720 5.380 ;
        RECT 82.420 5.030 84.720 5.270 ;
        RECT 82.420 4.930 82.870 5.030 ;
        RECT 83.260 4.600 83.670 5.030 ;
        RECT 84.270 4.960 84.720 5.030 ;
        RECT 85.670 5.270 86.120 5.350 ;
        RECT 86.720 5.270 87.130 5.710 ;
        RECT 87.520 5.270 87.970 5.380 ;
        RECT 85.670 5.030 87.970 5.270 ;
        RECT 85.670 4.930 86.120 5.030 ;
        RECT 87.520 4.930 87.970 5.030 ;
        RECT 89.160 5.270 89.610 5.380 ;
        RECT 90.000 5.270 90.410 5.710 ;
        RECT 93.180 5.440 93.630 5.720 ;
        RECT 97.000 5.440 97.450 5.720 ;
        RECT 106.680 5.720 108.210 5.930 ;
        RECT 108.590 5.840 109.040 5.930 ;
        RECT 109.420 5.720 110.950 5.930 ;
        RECT 91.010 5.270 91.460 5.350 ;
        RECT 89.160 5.030 91.460 5.270 ;
        RECT 89.160 4.930 89.610 5.030 ;
        RECT 91.010 4.930 91.460 5.030 ;
        RECT 92.410 5.270 92.860 5.380 ;
        RECT 94.260 5.270 94.710 5.380 ;
        RECT 92.410 5.030 94.710 5.270 ;
        RECT 92.410 4.960 92.860 5.030 ;
        RECT 75.660 4.400 76.110 4.450 ;
        RECT 74.020 4.110 76.110 4.400 ;
        RECT 74.020 4.060 74.470 4.110 ;
        RECT 57.270 3.480 57.720 3.550 ;
        RECT 55.420 3.240 57.720 3.480 ;
        RECT 55.420 3.130 55.870 3.240 ;
        RECT 57.270 3.130 57.720 3.240 ;
        RECT 58.670 3.480 59.120 3.580 ;
        RECT 60.520 3.480 60.970 3.580 ;
        RECT 58.670 3.240 60.970 3.480 ;
        RECT 58.670 3.160 59.120 3.240 ;
        RECT 39.180 2.580 40.710 2.790 ;
        RECT 41.090 2.580 41.540 2.670 ;
        RECT 41.920 2.580 43.450 2.790 ;
        RECT 52.680 2.790 53.130 3.070 ;
        RECT 56.500 2.790 56.950 3.070 ;
        RECT 59.720 2.800 60.130 3.240 ;
        RECT 60.520 3.130 60.970 3.240 ;
        RECT 62.160 3.480 62.610 3.580 ;
        RECT 64.010 3.480 64.460 3.580 ;
        RECT 62.160 3.240 64.460 3.480 ;
        RECT 62.160 3.130 62.610 3.240 ;
        RECT 63.000 2.800 63.410 3.240 ;
        RECT 64.010 3.160 64.460 3.240 ;
        RECT 65.410 3.480 65.860 3.550 ;
        RECT 66.460 3.480 66.870 3.910 ;
        RECT 67.260 3.480 67.710 3.580 ;
        RECT 65.410 3.240 67.710 3.480 ;
        RECT 65.410 3.130 65.860 3.240 ;
        RECT 67.260 3.130 67.710 3.240 ;
        RECT 68.920 3.480 69.370 3.580 ;
        RECT 69.760 3.480 70.170 3.910 ;
        RECT 72.920 3.840 74.470 4.060 ;
        RECT 74.850 4.050 75.280 4.110 ;
        RECT 75.660 4.060 76.110 4.110 ;
        RECT 76.710 4.060 77.210 4.450 ;
        RECT 75.660 3.840 77.210 4.060 ;
        RECT 86.420 4.450 87.970 4.670 ;
        RECT 86.420 4.060 86.920 4.450 ;
        RECT 87.520 4.400 87.970 4.450 ;
        RECT 88.350 4.400 88.780 4.460 ;
        RECT 89.160 4.450 90.710 4.670 ;
        RECT 93.460 4.600 93.870 5.030 ;
        RECT 94.260 4.930 94.710 5.030 ;
        RECT 95.920 5.270 96.370 5.380 ;
        RECT 97.770 5.270 98.220 5.380 ;
        RECT 95.920 5.030 98.220 5.270 ;
        RECT 95.920 4.930 96.370 5.030 ;
        RECT 96.760 4.600 97.170 5.030 ;
        RECT 97.770 4.960 98.220 5.030 ;
        RECT 99.170 5.270 99.620 5.350 ;
        RECT 100.220 5.270 100.630 5.710 ;
        RECT 101.020 5.270 101.470 5.380 ;
        RECT 99.170 5.030 101.470 5.270 ;
        RECT 99.170 4.930 99.620 5.030 ;
        RECT 101.020 4.930 101.470 5.030 ;
        RECT 102.660 5.270 103.110 5.380 ;
        RECT 103.500 5.270 103.910 5.710 ;
        RECT 106.680 5.440 107.130 5.720 ;
        RECT 110.500 5.440 110.950 5.720 ;
        RECT 120.180 5.720 121.710 5.930 ;
        RECT 122.090 5.840 122.540 5.930 ;
        RECT 122.920 5.720 124.450 5.930 ;
        RECT 104.510 5.270 104.960 5.350 ;
        RECT 102.660 5.030 104.960 5.270 ;
        RECT 102.660 4.930 103.110 5.030 ;
        RECT 104.510 4.930 104.960 5.030 ;
        RECT 105.910 5.270 106.360 5.380 ;
        RECT 107.760 5.270 108.210 5.380 ;
        RECT 105.910 5.030 108.210 5.270 ;
        RECT 105.910 4.960 106.360 5.030 ;
        RECT 89.160 4.400 89.610 4.450 ;
        RECT 87.520 4.110 89.610 4.400 ;
        RECT 87.520 4.060 87.970 4.110 ;
        RECT 70.770 3.480 71.220 3.550 ;
        RECT 68.920 3.240 71.220 3.480 ;
        RECT 68.920 3.130 69.370 3.240 ;
        RECT 70.770 3.130 71.220 3.240 ;
        RECT 72.170 3.480 72.620 3.580 ;
        RECT 74.020 3.480 74.470 3.580 ;
        RECT 72.170 3.240 74.470 3.480 ;
        RECT 72.170 3.160 72.620 3.240 ;
        RECT 52.680 2.630 54.210 2.790 ;
        RECT 54.590 2.630 55.040 2.670 ;
        RECT 55.420 2.630 56.950 2.790 ;
        RECT 52.680 2.580 56.950 2.630 ;
        RECT 66.180 2.790 66.630 3.070 ;
        RECT 70.000 2.790 70.450 3.070 ;
        RECT 73.220 2.800 73.630 3.240 ;
        RECT 74.020 3.130 74.470 3.240 ;
        RECT 75.660 3.480 76.110 3.580 ;
        RECT 77.510 3.480 77.960 3.580 ;
        RECT 75.660 3.240 77.960 3.480 ;
        RECT 75.660 3.130 76.110 3.240 ;
        RECT 76.500 2.800 76.910 3.240 ;
        RECT 77.510 3.160 77.960 3.240 ;
        RECT 78.910 3.480 79.360 3.550 ;
        RECT 79.960 3.480 80.370 3.910 ;
        RECT 80.760 3.480 81.210 3.580 ;
        RECT 78.910 3.240 81.210 3.480 ;
        RECT 78.910 3.130 79.360 3.240 ;
        RECT 80.760 3.130 81.210 3.240 ;
        RECT 82.420 3.480 82.870 3.580 ;
        RECT 83.260 3.480 83.670 3.910 ;
        RECT 86.420 3.840 87.970 4.060 ;
        RECT 88.350 4.050 88.780 4.110 ;
        RECT 89.160 4.060 89.610 4.110 ;
        RECT 90.210 4.060 90.710 4.450 ;
        RECT 89.160 3.840 90.710 4.060 ;
        RECT 99.920 4.450 101.470 4.670 ;
        RECT 99.920 4.060 100.420 4.450 ;
        RECT 101.020 4.400 101.470 4.450 ;
        RECT 101.850 4.400 102.280 4.460 ;
        RECT 102.660 4.450 104.210 4.670 ;
        RECT 106.960 4.600 107.370 5.030 ;
        RECT 107.760 4.930 108.210 5.030 ;
        RECT 109.420 5.270 109.870 5.380 ;
        RECT 111.270 5.270 111.720 5.380 ;
        RECT 109.420 5.030 111.720 5.270 ;
        RECT 109.420 4.930 109.870 5.030 ;
        RECT 110.260 4.600 110.670 5.030 ;
        RECT 111.270 4.960 111.720 5.030 ;
        RECT 112.670 5.270 113.120 5.350 ;
        RECT 113.720 5.270 114.130 5.710 ;
        RECT 114.520 5.270 114.970 5.380 ;
        RECT 112.670 5.030 114.970 5.270 ;
        RECT 112.670 4.930 113.120 5.030 ;
        RECT 114.520 4.930 114.970 5.030 ;
        RECT 116.160 5.270 116.610 5.380 ;
        RECT 117.000 5.270 117.410 5.710 ;
        RECT 120.180 5.440 120.630 5.720 ;
        RECT 124.000 5.440 124.450 5.720 ;
        RECT 133.680 5.720 135.210 5.930 ;
        RECT 135.590 5.840 136.040 5.930 ;
        RECT 136.420 5.720 137.950 5.930 ;
        RECT 118.010 5.270 118.460 5.350 ;
        RECT 116.160 5.030 118.460 5.270 ;
        RECT 116.160 4.930 116.610 5.030 ;
        RECT 118.010 4.930 118.460 5.030 ;
        RECT 119.410 5.270 119.860 5.380 ;
        RECT 121.260 5.270 121.710 5.380 ;
        RECT 119.410 5.030 121.710 5.270 ;
        RECT 119.410 4.960 119.860 5.030 ;
        RECT 102.660 4.400 103.110 4.450 ;
        RECT 101.020 4.110 103.110 4.400 ;
        RECT 101.020 4.060 101.470 4.110 ;
        RECT 84.270 3.480 84.720 3.550 ;
        RECT 82.420 3.240 84.720 3.480 ;
        RECT 82.420 3.130 82.870 3.240 ;
        RECT 84.270 3.130 84.720 3.240 ;
        RECT 85.670 3.480 86.120 3.580 ;
        RECT 87.520 3.480 87.970 3.580 ;
        RECT 85.670 3.240 87.970 3.480 ;
        RECT 85.670 3.160 86.120 3.240 ;
        RECT 66.180 2.580 67.710 2.790 ;
        RECT 68.090 2.580 68.540 2.670 ;
        RECT 68.920 2.580 70.450 2.790 ;
        RECT 79.680 2.790 80.130 3.070 ;
        RECT 83.500 2.790 83.950 3.070 ;
        RECT 86.720 2.800 87.130 3.240 ;
        RECT 87.520 3.130 87.970 3.240 ;
        RECT 89.160 3.480 89.610 3.580 ;
        RECT 91.010 3.480 91.460 3.580 ;
        RECT 89.160 3.240 91.460 3.480 ;
        RECT 89.160 3.130 89.610 3.240 ;
        RECT 90.000 2.800 90.410 3.240 ;
        RECT 91.010 3.160 91.460 3.240 ;
        RECT 92.410 3.480 92.860 3.550 ;
        RECT 93.460 3.480 93.870 3.910 ;
        RECT 94.260 3.480 94.710 3.580 ;
        RECT 92.410 3.240 94.710 3.480 ;
        RECT 92.410 3.130 92.860 3.240 ;
        RECT 94.260 3.130 94.710 3.240 ;
        RECT 95.920 3.480 96.370 3.580 ;
        RECT 96.760 3.480 97.170 3.910 ;
        RECT 99.920 3.840 101.470 4.060 ;
        RECT 101.850 4.050 102.280 4.110 ;
        RECT 102.660 4.060 103.110 4.110 ;
        RECT 103.710 4.060 104.210 4.450 ;
        RECT 102.660 3.840 104.210 4.060 ;
        RECT 113.420 4.450 114.970 4.670 ;
        RECT 113.420 4.060 113.920 4.450 ;
        RECT 114.520 4.400 114.970 4.450 ;
        RECT 115.350 4.400 115.780 4.460 ;
        RECT 116.160 4.450 117.710 4.670 ;
        RECT 120.460 4.600 120.870 5.030 ;
        RECT 121.260 4.930 121.710 5.030 ;
        RECT 122.920 5.270 123.370 5.380 ;
        RECT 124.770 5.270 125.220 5.380 ;
        RECT 122.920 5.030 125.220 5.270 ;
        RECT 122.920 4.930 123.370 5.030 ;
        RECT 123.760 4.600 124.170 5.030 ;
        RECT 124.770 4.960 125.220 5.030 ;
        RECT 126.170 5.270 126.620 5.350 ;
        RECT 127.220 5.270 127.630 5.710 ;
        RECT 128.020 5.270 128.470 5.380 ;
        RECT 126.170 5.030 128.470 5.270 ;
        RECT 126.170 4.930 126.620 5.030 ;
        RECT 128.020 4.930 128.470 5.030 ;
        RECT 129.660 5.270 130.110 5.380 ;
        RECT 130.500 5.270 130.910 5.710 ;
        RECT 133.680 5.440 134.130 5.720 ;
        RECT 137.500 5.440 137.950 5.720 ;
        RECT 147.180 5.720 148.710 5.930 ;
        RECT 149.090 5.840 149.540 5.930 ;
        RECT 149.920 5.720 151.450 5.930 ;
        RECT 131.510 5.270 131.960 5.350 ;
        RECT 129.660 5.030 131.960 5.270 ;
        RECT 129.660 4.930 130.110 5.030 ;
        RECT 131.510 4.930 131.960 5.030 ;
        RECT 132.910 5.270 133.360 5.380 ;
        RECT 134.760 5.270 135.210 5.380 ;
        RECT 132.910 5.030 135.210 5.270 ;
        RECT 132.910 4.960 133.360 5.030 ;
        RECT 116.160 4.400 116.610 4.450 ;
        RECT 114.520 4.110 116.610 4.400 ;
        RECT 114.520 4.060 114.970 4.110 ;
        RECT 97.770 3.480 98.220 3.550 ;
        RECT 95.920 3.240 98.220 3.480 ;
        RECT 95.920 3.130 96.370 3.240 ;
        RECT 97.770 3.130 98.220 3.240 ;
        RECT 99.170 3.480 99.620 3.580 ;
        RECT 101.020 3.480 101.470 3.580 ;
        RECT 99.170 3.240 101.470 3.480 ;
        RECT 99.170 3.160 99.620 3.240 ;
        RECT 79.680 2.580 81.210 2.790 ;
        RECT 81.590 2.580 82.040 2.670 ;
        RECT 82.420 2.580 83.950 2.790 ;
        RECT 93.180 2.790 93.630 3.070 ;
        RECT 97.000 2.790 97.450 3.070 ;
        RECT 100.220 2.800 100.630 3.240 ;
        RECT 101.020 3.130 101.470 3.240 ;
        RECT 102.660 3.480 103.110 3.580 ;
        RECT 104.510 3.480 104.960 3.580 ;
        RECT 102.660 3.240 104.960 3.480 ;
        RECT 102.660 3.130 103.110 3.240 ;
        RECT 103.500 2.800 103.910 3.240 ;
        RECT 104.510 3.160 104.960 3.240 ;
        RECT 105.910 3.480 106.360 3.550 ;
        RECT 106.960 3.480 107.370 3.910 ;
        RECT 107.760 3.480 108.210 3.580 ;
        RECT 105.910 3.240 108.210 3.480 ;
        RECT 105.910 3.130 106.360 3.240 ;
        RECT 107.760 3.130 108.210 3.240 ;
        RECT 109.420 3.480 109.870 3.580 ;
        RECT 110.260 3.480 110.670 3.910 ;
        RECT 113.420 3.840 114.970 4.060 ;
        RECT 115.350 4.050 115.780 4.110 ;
        RECT 116.160 4.060 116.610 4.110 ;
        RECT 117.210 4.060 117.710 4.450 ;
        RECT 116.160 3.840 117.710 4.060 ;
        RECT 126.920 4.450 128.470 4.670 ;
        RECT 126.920 4.060 127.420 4.450 ;
        RECT 128.020 4.400 128.470 4.450 ;
        RECT 128.850 4.400 129.280 4.460 ;
        RECT 129.660 4.450 131.210 4.670 ;
        RECT 133.960 4.600 134.370 5.030 ;
        RECT 134.760 4.930 135.210 5.030 ;
        RECT 136.420 5.270 136.870 5.380 ;
        RECT 138.270 5.270 138.720 5.380 ;
        RECT 136.420 5.030 138.720 5.270 ;
        RECT 136.420 4.930 136.870 5.030 ;
        RECT 137.260 4.600 137.670 5.030 ;
        RECT 138.270 4.960 138.720 5.030 ;
        RECT 139.670 5.270 140.120 5.350 ;
        RECT 140.720 5.270 141.130 5.710 ;
        RECT 141.520 5.270 141.970 5.380 ;
        RECT 139.670 5.030 141.970 5.270 ;
        RECT 139.670 4.930 140.120 5.030 ;
        RECT 141.520 4.930 141.970 5.030 ;
        RECT 143.160 5.270 143.610 5.380 ;
        RECT 144.000 5.270 144.410 5.710 ;
        RECT 147.180 5.440 147.630 5.720 ;
        RECT 151.000 5.440 151.450 5.720 ;
        RECT 160.680 5.720 162.210 5.930 ;
        RECT 162.590 5.840 163.040 5.930 ;
        RECT 163.420 5.720 164.950 5.930 ;
        RECT 145.010 5.270 145.460 5.350 ;
        RECT 143.160 5.030 145.460 5.270 ;
        RECT 143.160 4.930 143.610 5.030 ;
        RECT 145.010 4.930 145.460 5.030 ;
        RECT 146.410 5.270 146.860 5.380 ;
        RECT 148.260 5.270 148.710 5.380 ;
        RECT 146.410 5.030 148.710 5.270 ;
        RECT 146.410 4.960 146.860 5.030 ;
        RECT 129.660 4.400 130.110 4.450 ;
        RECT 128.020 4.110 130.110 4.400 ;
        RECT 128.020 4.060 128.470 4.110 ;
        RECT 111.270 3.480 111.720 3.550 ;
        RECT 109.420 3.240 111.720 3.480 ;
        RECT 109.420 3.130 109.870 3.240 ;
        RECT 111.270 3.130 111.720 3.240 ;
        RECT 112.670 3.480 113.120 3.580 ;
        RECT 114.520 3.480 114.970 3.580 ;
        RECT 112.670 3.240 114.970 3.480 ;
        RECT 112.670 3.160 113.120 3.240 ;
        RECT 93.180 2.580 94.710 2.790 ;
        RECT 95.090 2.580 95.540 2.670 ;
        RECT 95.920 2.580 97.450 2.790 ;
        RECT 106.680 2.790 107.130 3.070 ;
        RECT 110.500 2.790 110.950 3.070 ;
        RECT 113.720 2.800 114.130 3.240 ;
        RECT 114.520 3.130 114.970 3.240 ;
        RECT 116.160 3.480 116.610 3.580 ;
        RECT 118.010 3.480 118.460 3.580 ;
        RECT 116.160 3.240 118.460 3.480 ;
        RECT 116.160 3.130 116.610 3.240 ;
        RECT 117.000 2.800 117.410 3.240 ;
        RECT 118.010 3.160 118.460 3.240 ;
        RECT 119.410 3.480 119.860 3.550 ;
        RECT 120.460 3.480 120.870 3.910 ;
        RECT 121.260 3.480 121.710 3.580 ;
        RECT 119.410 3.240 121.710 3.480 ;
        RECT 119.410 3.130 119.860 3.240 ;
        RECT 121.260 3.130 121.710 3.240 ;
        RECT 122.920 3.480 123.370 3.580 ;
        RECT 123.760 3.480 124.170 3.910 ;
        RECT 126.920 3.840 128.470 4.060 ;
        RECT 128.850 4.050 129.280 4.110 ;
        RECT 129.660 4.060 130.110 4.110 ;
        RECT 130.710 4.060 131.210 4.450 ;
        RECT 129.660 3.840 131.210 4.060 ;
        RECT 140.420 4.450 141.970 4.670 ;
        RECT 140.420 4.060 140.920 4.450 ;
        RECT 141.520 4.400 141.970 4.450 ;
        RECT 142.350 4.400 142.780 4.460 ;
        RECT 143.160 4.450 144.710 4.670 ;
        RECT 147.460 4.600 147.870 5.030 ;
        RECT 148.260 4.930 148.710 5.030 ;
        RECT 149.920 5.270 150.370 5.380 ;
        RECT 151.770 5.270 152.220 5.380 ;
        RECT 149.920 5.030 152.220 5.270 ;
        RECT 149.920 4.930 150.370 5.030 ;
        RECT 150.760 4.600 151.170 5.030 ;
        RECT 151.770 4.960 152.220 5.030 ;
        RECT 153.170 5.270 153.620 5.350 ;
        RECT 154.220 5.270 154.630 5.710 ;
        RECT 155.020 5.270 155.470 5.380 ;
        RECT 153.170 5.030 155.470 5.270 ;
        RECT 153.170 4.930 153.620 5.030 ;
        RECT 155.020 4.930 155.470 5.030 ;
        RECT 156.660 5.270 157.110 5.380 ;
        RECT 157.500 5.270 157.910 5.710 ;
        RECT 160.680 5.440 161.130 5.720 ;
        RECT 164.500 5.440 164.950 5.720 ;
        RECT 174.180 5.720 175.710 5.930 ;
        RECT 176.090 5.840 176.540 5.930 ;
        RECT 176.920 5.720 178.450 5.930 ;
        RECT 158.510 5.270 158.960 5.350 ;
        RECT 156.660 5.030 158.960 5.270 ;
        RECT 156.660 4.930 157.110 5.030 ;
        RECT 158.510 4.930 158.960 5.030 ;
        RECT 159.910 5.270 160.360 5.380 ;
        RECT 161.760 5.270 162.210 5.380 ;
        RECT 159.910 5.030 162.210 5.270 ;
        RECT 159.910 4.960 160.360 5.030 ;
        RECT 143.160 4.400 143.610 4.450 ;
        RECT 141.520 4.110 143.610 4.400 ;
        RECT 141.520 4.060 141.970 4.110 ;
        RECT 124.770 3.480 125.220 3.550 ;
        RECT 122.920 3.240 125.220 3.480 ;
        RECT 122.920 3.130 123.370 3.240 ;
        RECT 124.770 3.130 125.220 3.240 ;
        RECT 126.170 3.480 126.620 3.580 ;
        RECT 128.020 3.480 128.470 3.580 ;
        RECT 126.170 3.240 128.470 3.480 ;
        RECT 126.170 3.160 126.620 3.240 ;
        RECT 106.680 2.630 108.210 2.790 ;
        RECT 108.590 2.630 109.040 2.670 ;
        RECT 109.420 2.630 110.950 2.790 ;
        RECT 106.680 2.580 110.950 2.630 ;
        RECT 120.180 2.790 120.630 3.070 ;
        RECT 124.000 2.790 124.450 3.070 ;
        RECT 127.220 2.800 127.630 3.240 ;
        RECT 128.020 3.130 128.470 3.240 ;
        RECT 129.660 3.480 130.110 3.580 ;
        RECT 131.510 3.480 131.960 3.580 ;
        RECT 129.660 3.240 131.960 3.480 ;
        RECT 129.660 3.130 130.110 3.240 ;
        RECT 130.500 2.800 130.910 3.240 ;
        RECT 131.510 3.160 131.960 3.240 ;
        RECT 132.910 3.480 133.360 3.550 ;
        RECT 133.960 3.480 134.370 3.910 ;
        RECT 134.760 3.480 135.210 3.580 ;
        RECT 132.910 3.240 135.210 3.480 ;
        RECT 132.910 3.130 133.360 3.240 ;
        RECT 134.760 3.130 135.210 3.240 ;
        RECT 136.420 3.480 136.870 3.580 ;
        RECT 137.260 3.480 137.670 3.910 ;
        RECT 140.420 3.840 141.970 4.060 ;
        RECT 142.350 4.050 142.780 4.110 ;
        RECT 143.160 4.060 143.610 4.110 ;
        RECT 144.210 4.060 144.710 4.450 ;
        RECT 143.160 3.840 144.710 4.060 ;
        RECT 153.920 4.450 155.470 4.670 ;
        RECT 153.920 4.060 154.420 4.450 ;
        RECT 155.020 4.400 155.470 4.450 ;
        RECT 155.850 4.400 156.280 4.460 ;
        RECT 156.660 4.450 158.210 4.670 ;
        RECT 160.960 4.600 161.370 5.030 ;
        RECT 161.760 4.930 162.210 5.030 ;
        RECT 163.420 5.270 163.870 5.380 ;
        RECT 165.270 5.270 165.720 5.380 ;
        RECT 163.420 5.030 165.720 5.270 ;
        RECT 163.420 4.930 163.870 5.030 ;
        RECT 164.260 4.600 164.670 5.030 ;
        RECT 165.270 4.960 165.720 5.030 ;
        RECT 166.670 5.270 167.120 5.350 ;
        RECT 167.720 5.270 168.130 5.710 ;
        RECT 168.520 5.270 168.970 5.380 ;
        RECT 166.670 5.030 168.970 5.270 ;
        RECT 166.670 4.930 167.120 5.030 ;
        RECT 168.520 4.930 168.970 5.030 ;
        RECT 170.160 5.270 170.610 5.380 ;
        RECT 171.000 5.270 171.410 5.710 ;
        RECT 174.180 5.440 174.630 5.720 ;
        RECT 178.000 5.440 178.450 5.720 ;
        RECT 187.680 5.720 189.210 5.930 ;
        RECT 189.590 5.840 190.040 5.930 ;
        RECT 190.420 5.720 191.950 5.930 ;
        RECT 172.010 5.270 172.460 5.350 ;
        RECT 170.160 5.030 172.460 5.270 ;
        RECT 170.160 4.930 170.610 5.030 ;
        RECT 172.010 4.930 172.460 5.030 ;
        RECT 173.410 5.270 173.860 5.380 ;
        RECT 175.260 5.270 175.710 5.380 ;
        RECT 173.410 5.030 175.710 5.270 ;
        RECT 173.410 4.960 173.860 5.030 ;
        RECT 156.660 4.400 157.110 4.450 ;
        RECT 155.020 4.110 157.110 4.400 ;
        RECT 155.020 4.060 155.470 4.110 ;
        RECT 138.270 3.480 138.720 3.550 ;
        RECT 136.420 3.240 138.720 3.480 ;
        RECT 136.420 3.130 136.870 3.240 ;
        RECT 138.270 3.130 138.720 3.240 ;
        RECT 139.670 3.480 140.120 3.580 ;
        RECT 141.520 3.480 141.970 3.580 ;
        RECT 139.670 3.240 141.970 3.480 ;
        RECT 139.670 3.160 140.120 3.240 ;
        RECT 120.180 2.580 121.710 2.790 ;
        RECT 122.090 2.580 122.540 2.670 ;
        RECT 122.920 2.580 124.450 2.790 ;
        RECT 133.680 2.790 134.130 3.070 ;
        RECT 137.500 2.790 137.950 3.070 ;
        RECT 140.720 2.800 141.130 3.240 ;
        RECT 141.520 3.130 141.970 3.240 ;
        RECT 143.160 3.480 143.610 3.580 ;
        RECT 145.010 3.480 145.460 3.580 ;
        RECT 143.160 3.240 145.460 3.480 ;
        RECT 143.160 3.130 143.610 3.240 ;
        RECT 144.000 2.800 144.410 3.240 ;
        RECT 145.010 3.160 145.460 3.240 ;
        RECT 146.410 3.480 146.860 3.550 ;
        RECT 147.460 3.480 147.870 3.910 ;
        RECT 148.260 3.480 148.710 3.580 ;
        RECT 146.410 3.240 148.710 3.480 ;
        RECT 146.410 3.130 146.860 3.240 ;
        RECT 148.260 3.130 148.710 3.240 ;
        RECT 149.920 3.480 150.370 3.580 ;
        RECT 150.760 3.480 151.170 3.910 ;
        RECT 153.920 3.840 155.470 4.060 ;
        RECT 155.850 4.050 156.280 4.110 ;
        RECT 156.660 4.060 157.110 4.110 ;
        RECT 157.710 4.060 158.210 4.450 ;
        RECT 156.660 3.840 158.210 4.060 ;
        RECT 167.420 4.450 168.970 4.670 ;
        RECT 167.420 4.060 167.920 4.450 ;
        RECT 168.520 4.400 168.970 4.450 ;
        RECT 169.350 4.400 169.780 4.460 ;
        RECT 170.160 4.450 171.710 4.670 ;
        RECT 174.460 4.600 174.870 5.030 ;
        RECT 175.260 4.930 175.710 5.030 ;
        RECT 176.920 5.270 177.370 5.380 ;
        RECT 178.770 5.270 179.220 5.380 ;
        RECT 176.920 5.030 179.220 5.270 ;
        RECT 176.920 4.930 177.370 5.030 ;
        RECT 177.760 4.600 178.170 5.030 ;
        RECT 178.770 4.960 179.220 5.030 ;
        RECT 180.170 5.270 180.620 5.350 ;
        RECT 181.220 5.270 181.630 5.710 ;
        RECT 182.020 5.270 182.470 5.380 ;
        RECT 180.170 5.030 182.470 5.270 ;
        RECT 180.170 4.930 180.620 5.030 ;
        RECT 182.020 4.930 182.470 5.030 ;
        RECT 183.660 5.270 184.110 5.380 ;
        RECT 184.500 5.270 184.910 5.710 ;
        RECT 187.680 5.440 188.130 5.720 ;
        RECT 191.500 5.440 191.950 5.720 ;
        RECT 201.180 5.720 202.710 5.930 ;
        RECT 203.090 5.840 203.540 5.930 ;
        RECT 203.920 5.720 205.450 5.930 ;
        RECT 185.510 5.270 185.960 5.350 ;
        RECT 183.660 5.030 185.960 5.270 ;
        RECT 183.660 4.930 184.110 5.030 ;
        RECT 185.510 4.930 185.960 5.030 ;
        RECT 186.910 5.270 187.360 5.380 ;
        RECT 188.760 5.270 189.210 5.380 ;
        RECT 186.910 5.030 189.210 5.270 ;
        RECT 186.910 4.960 187.360 5.030 ;
        RECT 170.160 4.400 170.610 4.450 ;
        RECT 168.520 4.110 170.610 4.400 ;
        RECT 168.520 4.060 168.970 4.110 ;
        RECT 151.770 3.480 152.220 3.550 ;
        RECT 149.920 3.240 152.220 3.480 ;
        RECT 149.920 3.130 150.370 3.240 ;
        RECT 151.770 3.130 152.220 3.240 ;
        RECT 153.170 3.480 153.620 3.580 ;
        RECT 155.020 3.480 155.470 3.580 ;
        RECT 153.170 3.240 155.470 3.480 ;
        RECT 153.170 3.160 153.620 3.240 ;
        RECT 133.680 2.580 135.210 2.790 ;
        RECT 135.590 2.580 136.040 2.670 ;
        RECT 136.420 2.580 137.950 2.790 ;
        RECT 147.180 2.790 147.630 3.070 ;
        RECT 151.000 2.790 151.450 3.070 ;
        RECT 154.220 2.800 154.630 3.240 ;
        RECT 155.020 3.130 155.470 3.240 ;
        RECT 156.660 3.480 157.110 3.580 ;
        RECT 158.510 3.480 158.960 3.580 ;
        RECT 156.660 3.240 158.960 3.480 ;
        RECT 156.660 3.130 157.110 3.240 ;
        RECT 157.500 2.800 157.910 3.240 ;
        RECT 158.510 3.160 158.960 3.240 ;
        RECT 159.910 3.480 160.360 3.550 ;
        RECT 160.960 3.480 161.370 3.910 ;
        RECT 161.760 3.480 162.210 3.580 ;
        RECT 159.910 3.240 162.210 3.480 ;
        RECT 159.910 3.130 160.360 3.240 ;
        RECT 161.760 3.130 162.210 3.240 ;
        RECT 163.420 3.480 163.870 3.580 ;
        RECT 164.260 3.480 164.670 3.910 ;
        RECT 167.420 3.840 168.970 4.060 ;
        RECT 169.350 4.050 169.780 4.110 ;
        RECT 170.160 4.060 170.610 4.110 ;
        RECT 171.210 4.060 171.710 4.450 ;
        RECT 170.160 3.840 171.710 4.060 ;
        RECT 180.920 4.450 182.470 4.670 ;
        RECT 180.920 4.060 181.420 4.450 ;
        RECT 182.020 4.400 182.470 4.450 ;
        RECT 182.850 4.400 183.280 4.460 ;
        RECT 183.660 4.450 185.210 4.670 ;
        RECT 187.960 4.600 188.370 5.030 ;
        RECT 188.760 4.930 189.210 5.030 ;
        RECT 190.420 5.270 190.870 5.380 ;
        RECT 192.270 5.270 192.720 5.380 ;
        RECT 190.420 5.030 192.720 5.270 ;
        RECT 190.420 4.930 190.870 5.030 ;
        RECT 191.260 4.600 191.670 5.030 ;
        RECT 192.270 4.960 192.720 5.030 ;
        RECT 193.670 5.270 194.120 5.350 ;
        RECT 194.720 5.270 195.130 5.710 ;
        RECT 195.520 5.270 195.970 5.380 ;
        RECT 193.670 5.030 195.970 5.270 ;
        RECT 193.670 4.930 194.120 5.030 ;
        RECT 195.520 4.930 195.970 5.030 ;
        RECT 197.160 5.270 197.610 5.380 ;
        RECT 198.000 5.270 198.410 5.710 ;
        RECT 201.180 5.440 201.630 5.720 ;
        RECT 205.000 5.440 205.450 5.720 ;
        RECT 214.680 5.720 216.210 5.930 ;
        RECT 216.590 5.840 217.030 5.930 ;
        RECT 199.010 5.270 199.460 5.350 ;
        RECT 197.160 5.030 199.460 5.270 ;
        RECT 197.160 4.930 197.610 5.030 ;
        RECT 199.010 4.930 199.460 5.030 ;
        RECT 200.410 5.270 200.860 5.380 ;
        RECT 202.260 5.270 202.710 5.380 ;
        RECT 200.410 5.030 202.710 5.270 ;
        RECT 200.410 4.960 200.860 5.030 ;
        RECT 183.660 4.400 184.110 4.450 ;
        RECT 182.020 4.110 184.110 4.400 ;
        RECT 182.020 4.060 182.470 4.110 ;
        RECT 165.270 3.480 165.720 3.550 ;
        RECT 163.420 3.240 165.720 3.480 ;
        RECT 163.420 3.130 163.870 3.240 ;
        RECT 165.270 3.130 165.720 3.240 ;
        RECT 166.670 3.480 167.120 3.580 ;
        RECT 168.520 3.480 168.970 3.580 ;
        RECT 166.670 3.240 168.970 3.480 ;
        RECT 166.670 3.160 167.120 3.240 ;
        RECT 147.180 2.580 148.710 2.790 ;
        RECT 149.090 2.580 149.540 2.670 ;
        RECT 149.920 2.580 151.450 2.790 ;
        RECT 160.680 2.790 161.130 3.070 ;
        RECT 164.500 2.790 164.950 3.070 ;
        RECT 167.720 2.800 168.130 3.240 ;
        RECT 168.520 3.130 168.970 3.240 ;
        RECT 170.160 3.480 170.610 3.580 ;
        RECT 172.010 3.480 172.460 3.580 ;
        RECT 170.160 3.240 172.460 3.480 ;
        RECT 170.160 3.130 170.610 3.240 ;
        RECT 171.000 2.800 171.410 3.240 ;
        RECT 172.010 3.160 172.460 3.240 ;
        RECT 173.410 3.480 173.860 3.550 ;
        RECT 174.460 3.480 174.870 3.910 ;
        RECT 175.260 3.480 175.710 3.580 ;
        RECT 173.410 3.240 175.710 3.480 ;
        RECT 173.410 3.130 173.860 3.240 ;
        RECT 175.260 3.130 175.710 3.240 ;
        RECT 176.920 3.480 177.370 3.580 ;
        RECT 177.760 3.480 178.170 3.910 ;
        RECT 180.920 3.840 182.470 4.060 ;
        RECT 182.850 4.050 183.280 4.110 ;
        RECT 183.660 4.060 184.110 4.110 ;
        RECT 184.710 4.060 185.210 4.450 ;
        RECT 183.660 3.840 185.210 4.060 ;
        RECT 194.420 4.450 195.970 4.670 ;
        RECT 194.420 4.060 194.920 4.450 ;
        RECT 195.520 4.400 195.970 4.450 ;
        RECT 196.350 4.400 196.780 4.460 ;
        RECT 197.160 4.450 198.710 4.670 ;
        RECT 201.460 4.600 201.870 5.030 ;
        RECT 202.260 4.930 202.710 5.030 ;
        RECT 203.920 5.270 204.370 5.380 ;
        RECT 205.770 5.270 206.220 5.380 ;
        RECT 203.920 5.030 206.220 5.270 ;
        RECT 203.920 4.930 204.370 5.030 ;
        RECT 204.760 4.600 205.170 5.030 ;
        RECT 205.770 4.960 206.220 5.030 ;
        RECT 207.170 5.270 207.620 5.350 ;
        RECT 208.220 5.270 208.630 5.710 ;
        RECT 209.020 5.270 209.470 5.380 ;
        RECT 207.170 5.030 209.470 5.270 ;
        RECT 207.170 4.930 207.620 5.030 ;
        RECT 209.020 4.930 209.470 5.030 ;
        RECT 210.660 5.270 211.110 5.380 ;
        RECT 211.500 5.270 211.910 5.710 ;
        RECT 214.680 5.440 215.130 5.720 ;
        RECT 212.510 5.270 212.960 5.350 ;
        RECT 210.660 5.030 212.960 5.270 ;
        RECT 210.660 4.930 211.110 5.030 ;
        RECT 212.510 4.930 212.960 5.030 ;
        RECT 213.910 5.270 214.360 5.380 ;
        RECT 215.760 5.270 216.210 5.380 ;
        RECT 213.910 5.030 216.210 5.270 ;
        RECT 213.910 4.960 214.360 5.030 ;
        RECT 197.160 4.400 197.610 4.450 ;
        RECT 195.520 4.110 197.610 4.400 ;
        RECT 195.520 4.060 195.970 4.110 ;
        RECT 178.770 3.480 179.220 3.550 ;
        RECT 176.920 3.240 179.220 3.480 ;
        RECT 176.920 3.130 177.370 3.240 ;
        RECT 178.770 3.130 179.220 3.240 ;
        RECT 180.170 3.480 180.620 3.580 ;
        RECT 182.020 3.480 182.470 3.580 ;
        RECT 180.170 3.240 182.470 3.480 ;
        RECT 180.170 3.160 180.620 3.240 ;
        RECT 160.680 2.630 162.210 2.790 ;
        RECT 162.590 2.630 163.040 2.670 ;
        RECT 163.420 2.630 164.950 2.790 ;
        RECT 160.680 2.580 164.950 2.630 ;
        RECT 174.180 2.790 174.630 3.070 ;
        RECT 178.000 2.790 178.450 3.070 ;
        RECT 181.220 2.800 181.630 3.240 ;
        RECT 182.020 3.130 182.470 3.240 ;
        RECT 183.660 3.480 184.110 3.580 ;
        RECT 185.510 3.480 185.960 3.580 ;
        RECT 183.660 3.240 185.960 3.480 ;
        RECT 183.660 3.130 184.110 3.240 ;
        RECT 184.500 2.800 184.910 3.240 ;
        RECT 185.510 3.160 185.960 3.240 ;
        RECT 186.910 3.480 187.360 3.550 ;
        RECT 187.960 3.480 188.370 3.910 ;
        RECT 188.760 3.480 189.210 3.580 ;
        RECT 186.910 3.240 189.210 3.480 ;
        RECT 186.910 3.130 187.360 3.240 ;
        RECT 188.760 3.130 189.210 3.240 ;
        RECT 190.420 3.480 190.870 3.580 ;
        RECT 191.260 3.480 191.670 3.910 ;
        RECT 194.420 3.840 195.970 4.060 ;
        RECT 196.350 4.050 196.780 4.110 ;
        RECT 197.160 4.060 197.610 4.110 ;
        RECT 198.210 4.060 198.710 4.450 ;
        RECT 197.160 3.840 198.710 4.060 ;
        RECT 207.920 4.450 209.470 4.670 ;
        RECT 207.920 4.060 208.420 4.450 ;
        RECT 209.020 4.400 209.470 4.450 ;
        RECT 209.850 4.400 210.280 4.460 ;
        RECT 210.660 4.450 212.210 4.670 ;
        RECT 214.960 4.600 215.370 5.030 ;
        RECT 215.760 4.930 216.210 5.030 ;
        RECT 210.660 4.400 211.110 4.450 ;
        RECT 209.020 4.110 211.110 4.400 ;
        RECT 209.020 4.060 209.470 4.110 ;
        RECT 192.270 3.480 192.720 3.550 ;
        RECT 190.420 3.240 192.720 3.480 ;
        RECT 190.420 3.130 190.870 3.240 ;
        RECT 192.270 3.130 192.720 3.240 ;
        RECT 193.670 3.480 194.120 3.580 ;
        RECT 195.520 3.480 195.970 3.580 ;
        RECT 193.670 3.240 195.970 3.480 ;
        RECT 193.670 3.160 194.120 3.240 ;
        RECT 174.180 2.580 175.710 2.790 ;
        RECT 176.090 2.580 176.540 2.670 ;
        RECT 176.920 2.580 178.450 2.790 ;
        RECT 187.680 2.790 188.130 3.070 ;
        RECT 191.500 2.790 191.950 3.070 ;
        RECT 194.720 2.800 195.130 3.240 ;
        RECT 195.520 3.130 195.970 3.240 ;
        RECT 197.160 3.480 197.610 3.580 ;
        RECT 199.010 3.480 199.460 3.580 ;
        RECT 197.160 3.240 199.460 3.480 ;
        RECT 197.160 3.130 197.610 3.240 ;
        RECT 198.000 2.800 198.410 3.240 ;
        RECT 199.010 3.160 199.460 3.240 ;
        RECT 200.410 3.480 200.860 3.550 ;
        RECT 201.460 3.480 201.870 3.910 ;
        RECT 202.260 3.480 202.710 3.580 ;
        RECT 200.410 3.240 202.710 3.480 ;
        RECT 200.410 3.130 200.860 3.240 ;
        RECT 202.260 3.130 202.710 3.240 ;
        RECT 203.920 3.480 204.370 3.580 ;
        RECT 204.760 3.480 205.170 3.910 ;
        RECT 207.920 3.840 209.470 4.060 ;
        RECT 209.850 4.050 210.280 4.110 ;
        RECT 210.660 4.060 211.110 4.110 ;
        RECT 211.710 4.060 212.210 4.450 ;
        RECT 210.660 3.840 212.210 4.060 ;
        RECT 205.770 3.480 206.220 3.550 ;
        RECT 203.920 3.240 206.220 3.480 ;
        RECT 203.920 3.130 204.370 3.240 ;
        RECT 205.770 3.130 206.220 3.240 ;
        RECT 207.170 3.480 207.620 3.580 ;
        RECT 209.020 3.480 209.470 3.580 ;
        RECT 207.170 3.240 209.470 3.480 ;
        RECT 207.170 3.160 207.620 3.240 ;
        RECT 187.680 2.580 189.210 2.790 ;
        RECT 189.590 2.580 190.040 2.670 ;
        RECT 190.420 2.580 191.950 2.790 ;
        RECT 201.180 2.790 201.630 3.070 ;
        RECT 205.000 2.790 205.450 3.070 ;
        RECT 208.220 2.800 208.630 3.240 ;
        RECT 209.020 3.130 209.470 3.240 ;
        RECT 210.660 3.480 211.110 3.580 ;
        RECT 212.510 3.480 212.960 3.580 ;
        RECT 210.660 3.240 212.960 3.480 ;
        RECT 210.660 3.130 211.110 3.240 ;
        RECT 211.500 2.800 211.910 3.240 ;
        RECT 212.510 3.160 212.960 3.240 ;
        RECT 213.910 3.480 214.360 3.550 ;
        RECT 214.960 3.480 215.370 3.910 ;
        RECT 215.760 3.480 216.210 3.580 ;
        RECT 213.910 3.240 216.210 3.480 ;
        RECT 213.910 3.130 214.360 3.240 ;
        RECT 215.760 3.130 216.210 3.240 ;
        RECT 201.180 2.580 202.710 2.790 ;
        RECT 203.090 2.580 203.540 2.670 ;
        RECT 203.920 2.580 205.450 2.790 ;
        RECT 214.680 2.790 215.130 3.070 ;
        RECT 214.680 2.580 216.210 2.790 ;
        RECT 216.590 2.630 217.030 2.670 ;
        RECT 216.590 2.580 217.690 2.630 ;
        RECT 13.260 2.320 15.370 2.580 ;
        RECT 26.760 2.320 28.870 2.580 ;
        RECT 40.260 2.320 42.370 2.580 ;
        RECT 53.760 2.320 55.870 2.580 ;
        RECT 67.260 2.320 69.370 2.580 ;
        RECT 80.760 2.320 82.870 2.580 ;
        RECT 94.260 2.320 96.370 2.580 ;
        RECT 107.760 2.320 109.870 2.580 ;
        RECT 121.260 2.320 123.370 2.580 ;
        RECT 134.760 2.320 136.870 2.580 ;
        RECT 148.260 2.320 150.370 2.580 ;
        RECT 161.760 2.320 163.870 2.580 ;
        RECT 175.260 2.320 177.370 2.580 ;
        RECT 188.760 2.320 190.870 2.580 ;
        RECT 202.260 2.320 204.370 2.580 ;
        RECT 215.760 2.320 217.690 2.580 ;
        RECT 12.180 2.110 13.710 2.320 ;
        RECT 14.090 2.230 14.540 2.320 ;
        RECT 14.920 2.110 16.450 2.320 ;
        RECT 1.420 1.660 1.870 1.770 ;
        RECT 3.270 1.660 3.720 1.770 ;
        RECT 1.420 1.420 3.720 1.660 ;
        RECT 1.420 1.320 1.870 1.420 ;
        RECT 2.260 0.990 2.670 1.420 ;
        RECT 3.270 1.350 3.720 1.420 ;
        RECT 4.670 1.660 5.120 1.740 ;
        RECT 5.720 1.660 6.130 2.100 ;
        RECT 6.520 1.660 6.970 1.770 ;
        RECT 4.670 1.420 6.970 1.660 ;
        RECT 4.670 1.320 5.120 1.420 ;
        RECT 6.520 1.320 6.970 1.420 ;
        RECT 8.160 1.660 8.610 1.770 ;
        RECT 9.000 1.660 9.410 2.100 ;
        RECT 12.180 1.830 12.630 2.110 ;
        RECT 16.000 1.830 16.450 2.110 ;
        RECT 25.680 2.110 27.210 2.320 ;
        RECT 27.590 2.230 28.040 2.320 ;
        RECT 28.420 2.110 29.950 2.320 ;
        RECT 10.010 1.660 10.460 1.740 ;
        RECT 8.160 1.420 10.460 1.660 ;
        RECT 8.160 1.320 8.610 1.420 ;
        RECT 10.010 1.320 10.460 1.420 ;
        RECT 11.410 1.660 11.860 1.770 ;
        RECT 13.260 1.660 13.710 1.770 ;
        RECT 11.410 1.420 13.710 1.660 ;
        RECT 11.410 1.350 11.860 1.420 ;
        RECT 5.420 0.840 6.970 1.060 ;
        RECT 5.420 0.450 5.920 0.840 ;
        RECT 6.520 0.790 6.970 0.840 ;
        RECT 7.350 0.790 7.780 0.850 ;
        RECT 8.160 0.840 9.710 1.060 ;
        RECT 12.460 0.990 12.870 1.420 ;
        RECT 13.260 1.320 13.710 1.420 ;
        RECT 14.920 1.660 15.370 1.770 ;
        RECT 16.770 1.660 17.220 1.770 ;
        RECT 14.920 1.420 17.220 1.660 ;
        RECT 14.920 1.320 15.370 1.420 ;
        RECT 15.760 0.990 16.170 1.420 ;
        RECT 16.770 1.350 17.220 1.420 ;
        RECT 18.170 1.660 18.620 1.740 ;
        RECT 19.220 1.660 19.630 2.100 ;
        RECT 20.020 1.660 20.470 1.770 ;
        RECT 18.170 1.420 20.470 1.660 ;
        RECT 18.170 1.320 18.620 1.420 ;
        RECT 20.020 1.320 20.470 1.420 ;
        RECT 21.660 1.660 22.110 1.770 ;
        RECT 22.500 1.660 22.910 2.100 ;
        RECT 25.680 1.830 26.130 2.110 ;
        RECT 29.500 1.830 29.950 2.110 ;
        RECT 39.180 2.110 40.710 2.320 ;
        RECT 41.090 2.230 41.540 2.320 ;
        RECT 41.920 2.110 43.450 2.320 ;
        RECT 23.510 1.660 23.960 1.740 ;
        RECT 21.660 1.420 23.960 1.660 ;
        RECT 21.660 1.320 22.110 1.420 ;
        RECT 23.510 1.320 23.960 1.420 ;
        RECT 24.910 1.660 25.360 1.770 ;
        RECT 26.760 1.660 27.210 1.770 ;
        RECT 24.910 1.420 27.210 1.660 ;
        RECT 24.910 1.350 25.360 1.420 ;
        RECT 8.160 0.790 8.610 0.840 ;
        RECT 6.520 0.500 8.610 0.790 ;
        RECT 6.520 0.450 6.970 0.500 ;
        RECT 1.420 -0.130 1.870 -0.030 ;
        RECT 2.260 -0.130 2.670 0.300 ;
        RECT 5.420 0.230 6.970 0.450 ;
        RECT 7.350 0.440 7.780 0.500 ;
        RECT 8.160 0.450 8.610 0.500 ;
        RECT 9.210 0.450 9.710 0.840 ;
        RECT 8.160 0.230 9.710 0.450 ;
        RECT 18.920 0.840 20.470 1.060 ;
        RECT 18.920 0.450 19.420 0.840 ;
        RECT 20.020 0.790 20.470 0.840 ;
        RECT 20.850 0.790 21.280 0.850 ;
        RECT 21.660 0.840 23.210 1.060 ;
        RECT 25.960 0.990 26.370 1.420 ;
        RECT 26.760 1.320 27.210 1.420 ;
        RECT 28.420 1.660 28.870 1.770 ;
        RECT 30.270 1.660 30.720 1.770 ;
        RECT 28.420 1.420 30.720 1.660 ;
        RECT 28.420 1.320 28.870 1.420 ;
        RECT 29.260 0.990 29.670 1.420 ;
        RECT 30.270 1.350 30.720 1.420 ;
        RECT 31.670 1.660 32.120 1.740 ;
        RECT 32.720 1.660 33.130 2.100 ;
        RECT 33.520 1.660 33.970 1.770 ;
        RECT 31.670 1.420 33.970 1.660 ;
        RECT 31.670 1.320 32.120 1.420 ;
        RECT 33.520 1.320 33.970 1.420 ;
        RECT 35.160 1.660 35.610 1.770 ;
        RECT 36.000 1.660 36.410 2.100 ;
        RECT 39.180 1.830 39.630 2.110 ;
        RECT 43.000 1.830 43.450 2.110 ;
        RECT 52.680 2.270 56.950 2.320 ;
        RECT 52.680 2.110 54.210 2.270 ;
        RECT 54.590 2.230 55.040 2.270 ;
        RECT 55.420 2.110 56.950 2.270 ;
        RECT 37.010 1.660 37.460 1.740 ;
        RECT 35.160 1.420 37.460 1.660 ;
        RECT 35.160 1.320 35.610 1.420 ;
        RECT 37.010 1.320 37.460 1.420 ;
        RECT 38.410 1.660 38.860 1.770 ;
        RECT 40.260 1.660 40.710 1.770 ;
        RECT 38.410 1.420 40.710 1.660 ;
        RECT 38.410 1.350 38.860 1.420 ;
        RECT 21.660 0.790 22.110 0.840 ;
        RECT 20.020 0.500 22.110 0.790 ;
        RECT 20.020 0.450 20.470 0.500 ;
        RECT 3.270 -0.130 3.720 -0.060 ;
        RECT 1.420 -0.370 3.720 -0.130 ;
        RECT 1.420 -0.480 1.870 -0.370 ;
        RECT 3.270 -0.480 3.720 -0.370 ;
        RECT 4.670 -0.130 5.120 -0.030 ;
        RECT 6.520 -0.130 6.970 -0.030 ;
        RECT 4.670 -0.370 6.970 -0.130 ;
        RECT 4.670 -0.450 5.120 -0.370 ;
        RECT 5.720 -0.810 6.130 -0.370 ;
        RECT 6.520 -0.480 6.970 -0.370 ;
        RECT 8.160 -0.130 8.610 -0.030 ;
        RECT 10.010 -0.130 10.460 -0.030 ;
        RECT 8.160 -0.370 10.460 -0.130 ;
        RECT 8.160 -0.480 8.610 -0.370 ;
        RECT 9.000 -0.810 9.410 -0.370 ;
        RECT 10.010 -0.450 10.460 -0.370 ;
        RECT 11.410 -0.130 11.860 -0.060 ;
        RECT 12.460 -0.130 12.870 0.300 ;
        RECT 13.260 -0.130 13.710 -0.030 ;
        RECT 11.410 -0.370 13.710 -0.130 ;
        RECT 11.410 -0.480 11.860 -0.370 ;
        RECT 13.260 -0.480 13.710 -0.370 ;
        RECT 14.920 -0.130 15.370 -0.030 ;
        RECT 15.760 -0.130 16.170 0.300 ;
        RECT 18.920 0.230 20.470 0.450 ;
        RECT 20.850 0.440 21.280 0.500 ;
        RECT 21.660 0.450 22.110 0.500 ;
        RECT 22.710 0.450 23.210 0.840 ;
        RECT 21.660 0.230 23.210 0.450 ;
        RECT 32.420 0.840 33.970 1.060 ;
        RECT 32.420 0.450 32.920 0.840 ;
        RECT 33.520 0.790 33.970 0.840 ;
        RECT 34.350 0.790 34.780 0.850 ;
        RECT 35.160 0.840 36.710 1.060 ;
        RECT 39.460 0.990 39.870 1.420 ;
        RECT 40.260 1.320 40.710 1.420 ;
        RECT 41.920 1.660 42.370 1.770 ;
        RECT 43.770 1.660 44.220 1.770 ;
        RECT 41.920 1.420 44.220 1.660 ;
        RECT 41.920 1.320 42.370 1.420 ;
        RECT 42.760 0.990 43.170 1.420 ;
        RECT 43.770 1.350 44.220 1.420 ;
        RECT 45.170 1.660 45.620 1.740 ;
        RECT 46.220 1.660 46.630 2.100 ;
        RECT 47.020 1.660 47.470 1.770 ;
        RECT 45.170 1.420 47.470 1.660 ;
        RECT 45.170 1.320 45.620 1.420 ;
        RECT 47.020 1.320 47.470 1.420 ;
        RECT 48.660 1.660 49.110 1.770 ;
        RECT 49.500 1.660 49.910 2.100 ;
        RECT 52.680 1.830 53.130 2.110 ;
        RECT 56.500 1.830 56.950 2.110 ;
        RECT 66.180 2.110 67.710 2.320 ;
        RECT 68.090 2.230 68.540 2.320 ;
        RECT 68.920 2.110 70.450 2.320 ;
        RECT 50.510 1.660 50.960 1.740 ;
        RECT 48.660 1.420 50.960 1.660 ;
        RECT 48.660 1.320 49.110 1.420 ;
        RECT 50.510 1.320 50.960 1.420 ;
        RECT 51.910 1.660 52.360 1.770 ;
        RECT 53.760 1.660 54.210 1.770 ;
        RECT 51.910 1.420 54.210 1.660 ;
        RECT 51.910 1.350 52.360 1.420 ;
        RECT 35.160 0.790 35.610 0.840 ;
        RECT 33.520 0.500 35.610 0.790 ;
        RECT 33.520 0.450 33.970 0.500 ;
        RECT 16.770 -0.130 17.220 -0.060 ;
        RECT 14.920 -0.370 17.220 -0.130 ;
        RECT 14.920 -0.480 15.370 -0.370 ;
        RECT 16.770 -0.480 17.220 -0.370 ;
        RECT 18.170 -0.130 18.620 -0.030 ;
        RECT 20.020 -0.130 20.470 -0.030 ;
        RECT 18.170 -0.370 20.470 -0.130 ;
        RECT 18.170 -0.450 18.620 -0.370 ;
        RECT 12.180 -0.820 12.630 -0.540 ;
        RECT 16.000 -0.820 16.450 -0.540 ;
        RECT 19.220 -0.810 19.630 -0.370 ;
        RECT 20.020 -0.480 20.470 -0.370 ;
        RECT 21.660 -0.130 22.110 -0.030 ;
        RECT 23.510 -0.130 23.960 -0.030 ;
        RECT 21.660 -0.370 23.960 -0.130 ;
        RECT 21.660 -0.480 22.110 -0.370 ;
        RECT 22.500 -0.810 22.910 -0.370 ;
        RECT 23.510 -0.450 23.960 -0.370 ;
        RECT 24.910 -0.130 25.360 -0.060 ;
        RECT 25.960 -0.130 26.370 0.300 ;
        RECT 26.760 -0.130 27.210 -0.030 ;
        RECT 24.910 -0.370 27.210 -0.130 ;
        RECT 24.910 -0.480 25.360 -0.370 ;
        RECT 26.760 -0.480 27.210 -0.370 ;
        RECT 28.420 -0.130 28.870 -0.030 ;
        RECT 29.260 -0.130 29.670 0.300 ;
        RECT 32.420 0.230 33.970 0.450 ;
        RECT 34.350 0.440 34.780 0.500 ;
        RECT 35.160 0.450 35.610 0.500 ;
        RECT 36.210 0.450 36.710 0.840 ;
        RECT 35.160 0.230 36.710 0.450 ;
        RECT 45.920 0.840 47.470 1.060 ;
        RECT 45.920 0.450 46.420 0.840 ;
        RECT 47.020 0.790 47.470 0.840 ;
        RECT 47.850 0.790 48.280 0.850 ;
        RECT 48.660 0.840 50.210 1.060 ;
        RECT 52.960 0.990 53.370 1.420 ;
        RECT 53.760 1.320 54.210 1.420 ;
        RECT 55.420 1.660 55.870 1.770 ;
        RECT 57.270 1.660 57.720 1.770 ;
        RECT 55.420 1.420 57.720 1.660 ;
        RECT 55.420 1.320 55.870 1.420 ;
        RECT 56.260 0.990 56.670 1.420 ;
        RECT 57.270 1.350 57.720 1.420 ;
        RECT 58.670 1.660 59.120 1.740 ;
        RECT 59.720 1.660 60.130 2.100 ;
        RECT 60.520 1.660 60.970 1.770 ;
        RECT 58.670 1.420 60.970 1.660 ;
        RECT 58.670 1.320 59.120 1.420 ;
        RECT 60.520 1.320 60.970 1.420 ;
        RECT 62.160 1.660 62.610 1.770 ;
        RECT 63.000 1.660 63.410 2.100 ;
        RECT 66.180 1.830 66.630 2.110 ;
        RECT 70.000 1.830 70.450 2.110 ;
        RECT 79.680 2.110 81.210 2.320 ;
        RECT 81.590 2.230 82.040 2.320 ;
        RECT 82.420 2.110 83.950 2.320 ;
        RECT 64.010 1.660 64.460 1.740 ;
        RECT 62.160 1.420 64.460 1.660 ;
        RECT 62.160 1.320 62.610 1.420 ;
        RECT 64.010 1.320 64.460 1.420 ;
        RECT 65.410 1.660 65.860 1.770 ;
        RECT 67.260 1.660 67.710 1.770 ;
        RECT 65.410 1.420 67.710 1.660 ;
        RECT 65.410 1.350 65.860 1.420 ;
        RECT 48.660 0.790 49.110 0.840 ;
        RECT 47.020 0.500 49.110 0.790 ;
        RECT 47.020 0.450 47.470 0.500 ;
        RECT 30.270 -0.130 30.720 -0.060 ;
        RECT 28.420 -0.370 30.720 -0.130 ;
        RECT 28.420 -0.480 28.870 -0.370 ;
        RECT 30.270 -0.480 30.720 -0.370 ;
        RECT 31.670 -0.130 32.120 -0.030 ;
        RECT 33.520 -0.130 33.970 -0.030 ;
        RECT 31.670 -0.370 33.970 -0.130 ;
        RECT 31.670 -0.450 32.120 -0.370 ;
        RECT 12.180 -1.030 13.710 -0.820 ;
        RECT 14.090 -1.030 14.540 -0.940 ;
        RECT 14.920 -1.030 16.450 -0.820 ;
        RECT 25.680 -0.820 26.130 -0.540 ;
        RECT 29.500 -0.820 29.950 -0.540 ;
        RECT 32.720 -0.810 33.130 -0.370 ;
        RECT 33.520 -0.480 33.970 -0.370 ;
        RECT 35.160 -0.130 35.610 -0.030 ;
        RECT 37.010 -0.130 37.460 -0.030 ;
        RECT 35.160 -0.370 37.460 -0.130 ;
        RECT 35.160 -0.480 35.610 -0.370 ;
        RECT 36.000 -0.810 36.410 -0.370 ;
        RECT 37.010 -0.450 37.460 -0.370 ;
        RECT 38.410 -0.130 38.860 -0.060 ;
        RECT 39.460 -0.130 39.870 0.300 ;
        RECT 40.260 -0.130 40.710 -0.030 ;
        RECT 38.410 -0.370 40.710 -0.130 ;
        RECT 38.410 -0.480 38.860 -0.370 ;
        RECT 40.260 -0.480 40.710 -0.370 ;
        RECT 41.920 -0.130 42.370 -0.030 ;
        RECT 42.760 -0.130 43.170 0.300 ;
        RECT 45.920 0.230 47.470 0.450 ;
        RECT 47.850 0.440 48.280 0.500 ;
        RECT 48.660 0.450 49.110 0.500 ;
        RECT 49.710 0.450 50.210 0.840 ;
        RECT 48.660 0.230 50.210 0.450 ;
        RECT 59.420 0.840 60.970 1.060 ;
        RECT 59.420 0.450 59.920 0.840 ;
        RECT 60.520 0.790 60.970 0.840 ;
        RECT 61.350 0.790 61.780 0.850 ;
        RECT 62.160 0.840 63.710 1.060 ;
        RECT 66.460 0.990 66.870 1.420 ;
        RECT 67.260 1.320 67.710 1.420 ;
        RECT 68.920 1.660 69.370 1.770 ;
        RECT 70.770 1.660 71.220 1.770 ;
        RECT 68.920 1.420 71.220 1.660 ;
        RECT 68.920 1.320 69.370 1.420 ;
        RECT 69.760 0.990 70.170 1.420 ;
        RECT 70.770 1.350 71.220 1.420 ;
        RECT 72.170 1.660 72.620 1.740 ;
        RECT 73.220 1.660 73.630 2.100 ;
        RECT 74.020 1.660 74.470 1.770 ;
        RECT 72.170 1.420 74.470 1.660 ;
        RECT 72.170 1.320 72.620 1.420 ;
        RECT 74.020 1.320 74.470 1.420 ;
        RECT 75.660 1.660 76.110 1.770 ;
        RECT 76.500 1.660 76.910 2.100 ;
        RECT 79.680 1.830 80.130 2.110 ;
        RECT 83.500 1.830 83.950 2.110 ;
        RECT 93.180 2.110 94.710 2.320 ;
        RECT 95.090 2.230 95.540 2.320 ;
        RECT 95.920 2.110 97.450 2.320 ;
        RECT 77.510 1.660 77.960 1.740 ;
        RECT 75.660 1.420 77.960 1.660 ;
        RECT 75.660 1.320 76.110 1.420 ;
        RECT 77.510 1.320 77.960 1.420 ;
        RECT 78.910 1.660 79.360 1.770 ;
        RECT 80.760 1.660 81.210 1.770 ;
        RECT 78.910 1.420 81.210 1.660 ;
        RECT 78.910 1.350 79.360 1.420 ;
        RECT 62.160 0.790 62.610 0.840 ;
        RECT 60.520 0.500 62.610 0.790 ;
        RECT 60.520 0.450 60.970 0.500 ;
        RECT 43.770 -0.130 44.220 -0.060 ;
        RECT 41.920 -0.370 44.220 -0.130 ;
        RECT 41.920 -0.480 42.370 -0.370 ;
        RECT 43.770 -0.480 44.220 -0.370 ;
        RECT 45.170 -0.130 45.620 -0.030 ;
        RECT 47.020 -0.130 47.470 -0.030 ;
        RECT 45.170 -0.370 47.470 -0.130 ;
        RECT 45.170 -0.450 45.620 -0.370 ;
        RECT 25.680 -1.030 27.210 -0.820 ;
        RECT 27.590 -1.030 28.040 -0.940 ;
        RECT 28.420 -1.030 29.950 -0.820 ;
        RECT 39.180 -0.820 39.630 -0.540 ;
        RECT 43.000 -0.820 43.450 -0.540 ;
        RECT 46.220 -0.810 46.630 -0.370 ;
        RECT 47.020 -0.480 47.470 -0.370 ;
        RECT 48.660 -0.130 49.110 -0.030 ;
        RECT 50.510 -0.130 50.960 -0.030 ;
        RECT 48.660 -0.370 50.960 -0.130 ;
        RECT 48.660 -0.480 49.110 -0.370 ;
        RECT 49.500 -0.810 49.910 -0.370 ;
        RECT 50.510 -0.450 50.960 -0.370 ;
        RECT 51.910 -0.130 52.360 -0.060 ;
        RECT 52.960 -0.130 53.370 0.300 ;
        RECT 53.760 -0.130 54.210 -0.030 ;
        RECT 51.910 -0.370 54.210 -0.130 ;
        RECT 51.910 -0.480 52.360 -0.370 ;
        RECT 53.760 -0.480 54.210 -0.370 ;
        RECT 55.420 -0.130 55.870 -0.030 ;
        RECT 56.260 -0.130 56.670 0.300 ;
        RECT 59.420 0.230 60.970 0.450 ;
        RECT 61.350 0.440 61.780 0.500 ;
        RECT 62.160 0.450 62.610 0.500 ;
        RECT 63.210 0.450 63.710 0.840 ;
        RECT 62.160 0.230 63.710 0.450 ;
        RECT 72.920 0.840 74.470 1.060 ;
        RECT 72.920 0.450 73.420 0.840 ;
        RECT 74.020 0.790 74.470 0.840 ;
        RECT 74.850 0.790 75.280 0.850 ;
        RECT 75.660 0.840 77.210 1.060 ;
        RECT 79.960 0.990 80.370 1.420 ;
        RECT 80.760 1.320 81.210 1.420 ;
        RECT 82.420 1.660 82.870 1.770 ;
        RECT 84.270 1.660 84.720 1.770 ;
        RECT 82.420 1.420 84.720 1.660 ;
        RECT 82.420 1.320 82.870 1.420 ;
        RECT 83.260 0.990 83.670 1.420 ;
        RECT 84.270 1.350 84.720 1.420 ;
        RECT 85.670 1.660 86.120 1.740 ;
        RECT 86.720 1.660 87.130 2.100 ;
        RECT 87.520 1.660 87.970 1.770 ;
        RECT 85.670 1.420 87.970 1.660 ;
        RECT 85.670 1.320 86.120 1.420 ;
        RECT 87.520 1.320 87.970 1.420 ;
        RECT 89.160 1.660 89.610 1.770 ;
        RECT 90.000 1.660 90.410 2.100 ;
        RECT 93.180 1.830 93.630 2.110 ;
        RECT 97.000 1.830 97.450 2.110 ;
        RECT 106.680 2.270 110.950 2.320 ;
        RECT 106.680 2.110 108.210 2.270 ;
        RECT 108.590 2.230 109.040 2.270 ;
        RECT 109.420 2.110 110.950 2.270 ;
        RECT 91.010 1.660 91.460 1.740 ;
        RECT 89.160 1.420 91.460 1.660 ;
        RECT 89.160 1.320 89.610 1.420 ;
        RECT 91.010 1.320 91.460 1.420 ;
        RECT 92.410 1.660 92.860 1.770 ;
        RECT 94.260 1.660 94.710 1.770 ;
        RECT 92.410 1.420 94.710 1.660 ;
        RECT 92.410 1.350 92.860 1.420 ;
        RECT 75.660 0.790 76.110 0.840 ;
        RECT 74.020 0.500 76.110 0.790 ;
        RECT 74.020 0.450 74.470 0.500 ;
        RECT 57.270 -0.130 57.720 -0.060 ;
        RECT 55.420 -0.370 57.720 -0.130 ;
        RECT 55.420 -0.480 55.870 -0.370 ;
        RECT 57.270 -0.480 57.720 -0.370 ;
        RECT 58.670 -0.130 59.120 -0.030 ;
        RECT 60.520 -0.130 60.970 -0.030 ;
        RECT 58.670 -0.370 60.970 -0.130 ;
        RECT 58.670 -0.450 59.120 -0.370 ;
        RECT 39.180 -1.030 40.710 -0.820 ;
        RECT 41.090 -1.030 41.540 -0.940 ;
        RECT 41.920 -1.030 43.450 -0.820 ;
        RECT 52.680 -0.820 53.130 -0.540 ;
        RECT 56.500 -0.820 56.950 -0.540 ;
        RECT 59.720 -0.810 60.130 -0.370 ;
        RECT 60.520 -0.480 60.970 -0.370 ;
        RECT 62.160 -0.130 62.610 -0.030 ;
        RECT 64.010 -0.130 64.460 -0.030 ;
        RECT 62.160 -0.370 64.460 -0.130 ;
        RECT 62.160 -0.480 62.610 -0.370 ;
        RECT 63.000 -0.810 63.410 -0.370 ;
        RECT 64.010 -0.450 64.460 -0.370 ;
        RECT 65.410 -0.130 65.860 -0.060 ;
        RECT 66.460 -0.130 66.870 0.300 ;
        RECT 67.260 -0.130 67.710 -0.030 ;
        RECT 65.410 -0.370 67.710 -0.130 ;
        RECT 65.410 -0.480 65.860 -0.370 ;
        RECT 67.260 -0.480 67.710 -0.370 ;
        RECT 68.920 -0.130 69.370 -0.030 ;
        RECT 69.760 -0.130 70.170 0.300 ;
        RECT 72.920 0.230 74.470 0.450 ;
        RECT 74.850 0.440 75.280 0.500 ;
        RECT 75.660 0.450 76.110 0.500 ;
        RECT 76.710 0.450 77.210 0.840 ;
        RECT 75.660 0.230 77.210 0.450 ;
        RECT 86.420 0.840 87.970 1.060 ;
        RECT 86.420 0.450 86.920 0.840 ;
        RECT 87.520 0.790 87.970 0.840 ;
        RECT 88.350 0.790 88.780 0.850 ;
        RECT 89.160 0.840 90.710 1.060 ;
        RECT 93.460 0.990 93.870 1.420 ;
        RECT 94.260 1.320 94.710 1.420 ;
        RECT 95.920 1.660 96.370 1.770 ;
        RECT 97.770 1.660 98.220 1.770 ;
        RECT 95.920 1.420 98.220 1.660 ;
        RECT 95.920 1.320 96.370 1.420 ;
        RECT 96.760 0.990 97.170 1.420 ;
        RECT 97.770 1.350 98.220 1.420 ;
        RECT 99.170 1.660 99.620 1.740 ;
        RECT 100.220 1.660 100.630 2.100 ;
        RECT 101.020 1.660 101.470 1.770 ;
        RECT 99.170 1.420 101.470 1.660 ;
        RECT 99.170 1.320 99.620 1.420 ;
        RECT 101.020 1.320 101.470 1.420 ;
        RECT 102.660 1.660 103.110 1.770 ;
        RECT 103.500 1.660 103.910 2.100 ;
        RECT 106.680 1.830 107.130 2.110 ;
        RECT 110.500 1.830 110.950 2.110 ;
        RECT 120.180 2.110 121.710 2.320 ;
        RECT 122.090 2.230 122.540 2.320 ;
        RECT 122.920 2.110 124.450 2.320 ;
        RECT 104.510 1.660 104.960 1.740 ;
        RECT 102.660 1.420 104.960 1.660 ;
        RECT 102.660 1.320 103.110 1.420 ;
        RECT 104.510 1.320 104.960 1.420 ;
        RECT 105.910 1.660 106.360 1.770 ;
        RECT 107.760 1.660 108.210 1.770 ;
        RECT 105.910 1.420 108.210 1.660 ;
        RECT 105.910 1.350 106.360 1.420 ;
        RECT 89.160 0.790 89.610 0.840 ;
        RECT 87.520 0.500 89.610 0.790 ;
        RECT 87.520 0.450 87.970 0.500 ;
        RECT 70.770 -0.130 71.220 -0.060 ;
        RECT 68.920 -0.370 71.220 -0.130 ;
        RECT 68.920 -0.480 69.370 -0.370 ;
        RECT 70.770 -0.480 71.220 -0.370 ;
        RECT 72.170 -0.130 72.620 -0.030 ;
        RECT 74.020 -0.130 74.470 -0.030 ;
        RECT 72.170 -0.370 74.470 -0.130 ;
        RECT 72.170 -0.450 72.620 -0.370 ;
        RECT 52.680 -1.030 54.210 -0.820 ;
        RECT 54.590 -1.030 55.040 -0.940 ;
        RECT 55.420 -1.030 56.950 -0.820 ;
        RECT 66.180 -0.820 66.630 -0.540 ;
        RECT 70.000 -0.820 70.450 -0.540 ;
        RECT 73.220 -0.810 73.630 -0.370 ;
        RECT 74.020 -0.480 74.470 -0.370 ;
        RECT 75.660 -0.130 76.110 -0.030 ;
        RECT 77.510 -0.130 77.960 -0.030 ;
        RECT 75.660 -0.370 77.960 -0.130 ;
        RECT 75.660 -0.480 76.110 -0.370 ;
        RECT 76.500 -0.810 76.910 -0.370 ;
        RECT 77.510 -0.450 77.960 -0.370 ;
        RECT 78.910 -0.130 79.360 -0.060 ;
        RECT 79.960 -0.130 80.370 0.300 ;
        RECT 80.760 -0.130 81.210 -0.030 ;
        RECT 78.910 -0.370 81.210 -0.130 ;
        RECT 78.910 -0.480 79.360 -0.370 ;
        RECT 80.760 -0.480 81.210 -0.370 ;
        RECT 82.420 -0.130 82.870 -0.030 ;
        RECT 83.260 -0.130 83.670 0.300 ;
        RECT 86.420 0.230 87.970 0.450 ;
        RECT 88.350 0.440 88.780 0.500 ;
        RECT 89.160 0.450 89.610 0.500 ;
        RECT 90.210 0.450 90.710 0.840 ;
        RECT 89.160 0.230 90.710 0.450 ;
        RECT 99.920 0.840 101.470 1.060 ;
        RECT 99.920 0.450 100.420 0.840 ;
        RECT 101.020 0.790 101.470 0.840 ;
        RECT 101.850 0.790 102.280 0.850 ;
        RECT 102.660 0.840 104.210 1.060 ;
        RECT 106.960 0.990 107.370 1.420 ;
        RECT 107.760 1.320 108.210 1.420 ;
        RECT 109.420 1.660 109.870 1.770 ;
        RECT 111.270 1.660 111.720 1.770 ;
        RECT 109.420 1.420 111.720 1.660 ;
        RECT 109.420 1.320 109.870 1.420 ;
        RECT 110.260 0.990 110.670 1.420 ;
        RECT 111.270 1.350 111.720 1.420 ;
        RECT 112.670 1.660 113.120 1.740 ;
        RECT 113.720 1.660 114.130 2.100 ;
        RECT 114.520 1.660 114.970 1.770 ;
        RECT 112.670 1.420 114.970 1.660 ;
        RECT 112.670 1.320 113.120 1.420 ;
        RECT 114.520 1.320 114.970 1.420 ;
        RECT 116.160 1.660 116.610 1.770 ;
        RECT 117.000 1.660 117.410 2.100 ;
        RECT 120.180 1.830 120.630 2.110 ;
        RECT 124.000 1.830 124.450 2.110 ;
        RECT 133.680 2.110 135.210 2.320 ;
        RECT 135.590 2.230 136.040 2.320 ;
        RECT 136.420 2.110 137.950 2.320 ;
        RECT 118.010 1.660 118.460 1.740 ;
        RECT 116.160 1.420 118.460 1.660 ;
        RECT 116.160 1.320 116.610 1.420 ;
        RECT 118.010 1.320 118.460 1.420 ;
        RECT 119.410 1.660 119.860 1.770 ;
        RECT 121.260 1.660 121.710 1.770 ;
        RECT 119.410 1.420 121.710 1.660 ;
        RECT 119.410 1.350 119.860 1.420 ;
        RECT 102.660 0.790 103.110 0.840 ;
        RECT 101.020 0.500 103.110 0.790 ;
        RECT 101.020 0.450 101.470 0.500 ;
        RECT 84.270 -0.130 84.720 -0.060 ;
        RECT 82.420 -0.370 84.720 -0.130 ;
        RECT 82.420 -0.480 82.870 -0.370 ;
        RECT 84.270 -0.480 84.720 -0.370 ;
        RECT 85.670 -0.130 86.120 -0.030 ;
        RECT 87.520 -0.130 87.970 -0.030 ;
        RECT 85.670 -0.370 87.970 -0.130 ;
        RECT 85.670 -0.450 86.120 -0.370 ;
        RECT 66.180 -1.030 67.710 -0.820 ;
        RECT 68.090 -1.030 68.540 -0.940 ;
        RECT 68.920 -1.030 70.450 -0.820 ;
        RECT 79.680 -0.820 80.130 -0.540 ;
        RECT 83.500 -0.820 83.950 -0.540 ;
        RECT 86.720 -0.810 87.130 -0.370 ;
        RECT 87.520 -0.480 87.970 -0.370 ;
        RECT 89.160 -0.130 89.610 -0.030 ;
        RECT 91.010 -0.130 91.460 -0.030 ;
        RECT 89.160 -0.370 91.460 -0.130 ;
        RECT 89.160 -0.480 89.610 -0.370 ;
        RECT 90.000 -0.810 90.410 -0.370 ;
        RECT 91.010 -0.450 91.460 -0.370 ;
        RECT 92.410 -0.130 92.860 -0.060 ;
        RECT 93.460 -0.130 93.870 0.300 ;
        RECT 94.260 -0.130 94.710 -0.030 ;
        RECT 92.410 -0.370 94.710 -0.130 ;
        RECT 92.410 -0.480 92.860 -0.370 ;
        RECT 94.260 -0.480 94.710 -0.370 ;
        RECT 95.920 -0.130 96.370 -0.030 ;
        RECT 96.760 -0.130 97.170 0.300 ;
        RECT 99.920 0.230 101.470 0.450 ;
        RECT 101.850 0.440 102.280 0.500 ;
        RECT 102.660 0.450 103.110 0.500 ;
        RECT 103.710 0.450 104.210 0.840 ;
        RECT 102.660 0.230 104.210 0.450 ;
        RECT 113.420 0.840 114.970 1.060 ;
        RECT 113.420 0.450 113.920 0.840 ;
        RECT 114.520 0.790 114.970 0.840 ;
        RECT 115.350 0.790 115.780 0.850 ;
        RECT 116.160 0.840 117.710 1.060 ;
        RECT 120.460 0.990 120.870 1.420 ;
        RECT 121.260 1.320 121.710 1.420 ;
        RECT 122.920 1.660 123.370 1.770 ;
        RECT 124.770 1.660 125.220 1.770 ;
        RECT 122.920 1.420 125.220 1.660 ;
        RECT 122.920 1.320 123.370 1.420 ;
        RECT 123.760 0.990 124.170 1.420 ;
        RECT 124.770 1.350 125.220 1.420 ;
        RECT 126.170 1.660 126.620 1.740 ;
        RECT 127.220 1.660 127.630 2.100 ;
        RECT 128.020 1.660 128.470 1.770 ;
        RECT 126.170 1.420 128.470 1.660 ;
        RECT 126.170 1.320 126.620 1.420 ;
        RECT 128.020 1.320 128.470 1.420 ;
        RECT 129.660 1.660 130.110 1.770 ;
        RECT 130.500 1.660 130.910 2.100 ;
        RECT 133.680 1.830 134.130 2.110 ;
        RECT 137.500 1.830 137.950 2.110 ;
        RECT 147.180 2.110 148.710 2.320 ;
        RECT 149.090 2.230 149.540 2.320 ;
        RECT 149.920 2.110 151.450 2.320 ;
        RECT 131.510 1.660 131.960 1.740 ;
        RECT 129.660 1.420 131.960 1.660 ;
        RECT 129.660 1.320 130.110 1.420 ;
        RECT 131.510 1.320 131.960 1.420 ;
        RECT 132.910 1.660 133.360 1.770 ;
        RECT 134.760 1.660 135.210 1.770 ;
        RECT 132.910 1.420 135.210 1.660 ;
        RECT 132.910 1.350 133.360 1.420 ;
        RECT 116.160 0.790 116.610 0.840 ;
        RECT 114.520 0.500 116.610 0.790 ;
        RECT 114.520 0.450 114.970 0.500 ;
        RECT 97.770 -0.130 98.220 -0.060 ;
        RECT 95.920 -0.370 98.220 -0.130 ;
        RECT 95.920 -0.480 96.370 -0.370 ;
        RECT 97.770 -0.480 98.220 -0.370 ;
        RECT 99.170 -0.130 99.620 -0.030 ;
        RECT 101.020 -0.130 101.470 -0.030 ;
        RECT 99.170 -0.370 101.470 -0.130 ;
        RECT 99.170 -0.450 99.620 -0.370 ;
        RECT 79.680 -1.030 81.210 -0.820 ;
        RECT 81.590 -1.030 82.040 -0.940 ;
        RECT 82.420 -1.030 83.950 -0.820 ;
        RECT 93.180 -0.820 93.630 -0.540 ;
        RECT 97.000 -0.820 97.450 -0.540 ;
        RECT 100.220 -0.810 100.630 -0.370 ;
        RECT 101.020 -0.480 101.470 -0.370 ;
        RECT 102.660 -0.130 103.110 -0.030 ;
        RECT 104.510 -0.130 104.960 -0.030 ;
        RECT 102.660 -0.370 104.960 -0.130 ;
        RECT 102.660 -0.480 103.110 -0.370 ;
        RECT 103.500 -0.810 103.910 -0.370 ;
        RECT 104.510 -0.450 104.960 -0.370 ;
        RECT 105.910 -0.130 106.360 -0.060 ;
        RECT 106.960 -0.130 107.370 0.300 ;
        RECT 107.760 -0.130 108.210 -0.030 ;
        RECT 105.910 -0.370 108.210 -0.130 ;
        RECT 105.910 -0.480 106.360 -0.370 ;
        RECT 107.760 -0.480 108.210 -0.370 ;
        RECT 109.420 -0.130 109.870 -0.030 ;
        RECT 110.260 -0.130 110.670 0.300 ;
        RECT 113.420 0.230 114.970 0.450 ;
        RECT 115.350 0.440 115.780 0.500 ;
        RECT 116.160 0.450 116.610 0.500 ;
        RECT 117.210 0.450 117.710 0.840 ;
        RECT 116.160 0.230 117.710 0.450 ;
        RECT 126.920 0.840 128.470 1.060 ;
        RECT 126.920 0.450 127.420 0.840 ;
        RECT 128.020 0.790 128.470 0.840 ;
        RECT 128.850 0.790 129.280 0.850 ;
        RECT 129.660 0.840 131.210 1.060 ;
        RECT 133.960 0.990 134.370 1.420 ;
        RECT 134.760 1.320 135.210 1.420 ;
        RECT 136.420 1.660 136.870 1.770 ;
        RECT 138.270 1.660 138.720 1.770 ;
        RECT 136.420 1.420 138.720 1.660 ;
        RECT 136.420 1.320 136.870 1.420 ;
        RECT 137.260 0.990 137.670 1.420 ;
        RECT 138.270 1.350 138.720 1.420 ;
        RECT 139.670 1.660 140.120 1.740 ;
        RECT 140.720 1.660 141.130 2.100 ;
        RECT 141.520 1.660 141.970 1.770 ;
        RECT 139.670 1.420 141.970 1.660 ;
        RECT 139.670 1.320 140.120 1.420 ;
        RECT 141.520 1.320 141.970 1.420 ;
        RECT 143.160 1.660 143.610 1.770 ;
        RECT 144.000 1.660 144.410 2.100 ;
        RECT 147.180 1.830 147.630 2.110 ;
        RECT 151.000 1.830 151.450 2.110 ;
        RECT 160.680 2.270 164.950 2.320 ;
        RECT 160.680 2.110 162.210 2.270 ;
        RECT 162.590 2.230 163.040 2.270 ;
        RECT 163.420 2.110 164.950 2.270 ;
        RECT 145.010 1.660 145.460 1.740 ;
        RECT 143.160 1.420 145.460 1.660 ;
        RECT 143.160 1.320 143.610 1.420 ;
        RECT 145.010 1.320 145.460 1.420 ;
        RECT 146.410 1.660 146.860 1.770 ;
        RECT 148.260 1.660 148.710 1.770 ;
        RECT 146.410 1.420 148.710 1.660 ;
        RECT 146.410 1.350 146.860 1.420 ;
        RECT 129.660 0.790 130.110 0.840 ;
        RECT 128.020 0.500 130.110 0.790 ;
        RECT 128.020 0.450 128.470 0.500 ;
        RECT 111.270 -0.130 111.720 -0.060 ;
        RECT 109.420 -0.370 111.720 -0.130 ;
        RECT 109.420 -0.480 109.870 -0.370 ;
        RECT 111.270 -0.480 111.720 -0.370 ;
        RECT 112.670 -0.130 113.120 -0.030 ;
        RECT 114.520 -0.130 114.970 -0.030 ;
        RECT 112.670 -0.370 114.970 -0.130 ;
        RECT 112.670 -0.450 113.120 -0.370 ;
        RECT 93.180 -1.030 94.710 -0.820 ;
        RECT 95.090 -1.030 95.540 -0.940 ;
        RECT 95.920 -1.030 97.450 -0.820 ;
        RECT 106.680 -0.820 107.130 -0.540 ;
        RECT 110.500 -0.820 110.950 -0.540 ;
        RECT 113.720 -0.810 114.130 -0.370 ;
        RECT 114.520 -0.480 114.970 -0.370 ;
        RECT 116.160 -0.130 116.610 -0.030 ;
        RECT 118.010 -0.130 118.460 -0.030 ;
        RECT 116.160 -0.370 118.460 -0.130 ;
        RECT 116.160 -0.480 116.610 -0.370 ;
        RECT 117.000 -0.810 117.410 -0.370 ;
        RECT 118.010 -0.450 118.460 -0.370 ;
        RECT 119.410 -0.130 119.860 -0.060 ;
        RECT 120.460 -0.130 120.870 0.300 ;
        RECT 121.260 -0.130 121.710 -0.030 ;
        RECT 119.410 -0.370 121.710 -0.130 ;
        RECT 119.410 -0.480 119.860 -0.370 ;
        RECT 121.260 -0.480 121.710 -0.370 ;
        RECT 122.920 -0.130 123.370 -0.030 ;
        RECT 123.760 -0.130 124.170 0.300 ;
        RECT 126.920 0.230 128.470 0.450 ;
        RECT 128.850 0.440 129.280 0.500 ;
        RECT 129.660 0.450 130.110 0.500 ;
        RECT 130.710 0.450 131.210 0.840 ;
        RECT 129.660 0.230 131.210 0.450 ;
        RECT 140.420 0.840 141.970 1.060 ;
        RECT 140.420 0.450 140.920 0.840 ;
        RECT 141.520 0.790 141.970 0.840 ;
        RECT 142.350 0.790 142.780 0.850 ;
        RECT 143.160 0.840 144.710 1.060 ;
        RECT 147.460 0.990 147.870 1.420 ;
        RECT 148.260 1.320 148.710 1.420 ;
        RECT 149.920 1.660 150.370 1.770 ;
        RECT 151.770 1.660 152.220 1.770 ;
        RECT 149.920 1.420 152.220 1.660 ;
        RECT 149.920 1.320 150.370 1.420 ;
        RECT 150.760 0.990 151.170 1.420 ;
        RECT 151.770 1.350 152.220 1.420 ;
        RECT 153.170 1.660 153.620 1.740 ;
        RECT 154.220 1.660 154.630 2.100 ;
        RECT 155.020 1.660 155.470 1.770 ;
        RECT 153.170 1.420 155.470 1.660 ;
        RECT 153.170 1.320 153.620 1.420 ;
        RECT 155.020 1.320 155.470 1.420 ;
        RECT 156.660 1.660 157.110 1.770 ;
        RECT 157.500 1.660 157.910 2.100 ;
        RECT 160.680 1.830 161.130 2.110 ;
        RECT 164.500 1.830 164.950 2.110 ;
        RECT 174.180 2.110 175.710 2.320 ;
        RECT 176.090 2.230 176.540 2.320 ;
        RECT 176.920 2.110 178.450 2.320 ;
        RECT 158.510 1.660 158.960 1.740 ;
        RECT 156.660 1.420 158.960 1.660 ;
        RECT 156.660 1.320 157.110 1.420 ;
        RECT 158.510 1.320 158.960 1.420 ;
        RECT 159.910 1.660 160.360 1.770 ;
        RECT 161.760 1.660 162.210 1.770 ;
        RECT 159.910 1.420 162.210 1.660 ;
        RECT 159.910 1.350 160.360 1.420 ;
        RECT 143.160 0.790 143.610 0.840 ;
        RECT 141.520 0.500 143.610 0.790 ;
        RECT 141.520 0.450 141.970 0.500 ;
        RECT 124.770 -0.130 125.220 -0.060 ;
        RECT 122.920 -0.370 125.220 -0.130 ;
        RECT 122.920 -0.480 123.370 -0.370 ;
        RECT 124.770 -0.480 125.220 -0.370 ;
        RECT 126.170 -0.130 126.620 -0.030 ;
        RECT 128.020 -0.130 128.470 -0.030 ;
        RECT 126.170 -0.370 128.470 -0.130 ;
        RECT 126.170 -0.450 126.620 -0.370 ;
        RECT 106.680 -1.030 108.210 -0.820 ;
        RECT 108.590 -1.030 109.040 -0.940 ;
        RECT 109.420 -1.030 110.950 -0.820 ;
        RECT 120.180 -0.820 120.630 -0.540 ;
        RECT 124.000 -0.820 124.450 -0.540 ;
        RECT 127.220 -0.810 127.630 -0.370 ;
        RECT 128.020 -0.480 128.470 -0.370 ;
        RECT 129.660 -0.130 130.110 -0.030 ;
        RECT 131.510 -0.130 131.960 -0.030 ;
        RECT 129.660 -0.370 131.960 -0.130 ;
        RECT 129.660 -0.480 130.110 -0.370 ;
        RECT 130.500 -0.810 130.910 -0.370 ;
        RECT 131.510 -0.450 131.960 -0.370 ;
        RECT 132.910 -0.130 133.360 -0.060 ;
        RECT 133.960 -0.130 134.370 0.300 ;
        RECT 134.760 -0.130 135.210 -0.030 ;
        RECT 132.910 -0.370 135.210 -0.130 ;
        RECT 132.910 -0.480 133.360 -0.370 ;
        RECT 134.760 -0.480 135.210 -0.370 ;
        RECT 136.420 -0.130 136.870 -0.030 ;
        RECT 137.260 -0.130 137.670 0.300 ;
        RECT 140.420 0.230 141.970 0.450 ;
        RECT 142.350 0.440 142.780 0.500 ;
        RECT 143.160 0.450 143.610 0.500 ;
        RECT 144.210 0.450 144.710 0.840 ;
        RECT 143.160 0.230 144.710 0.450 ;
        RECT 153.920 0.840 155.470 1.060 ;
        RECT 153.920 0.450 154.420 0.840 ;
        RECT 155.020 0.790 155.470 0.840 ;
        RECT 155.850 0.790 156.280 0.850 ;
        RECT 156.660 0.840 158.210 1.060 ;
        RECT 160.960 0.990 161.370 1.420 ;
        RECT 161.760 1.320 162.210 1.420 ;
        RECT 163.420 1.660 163.870 1.770 ;
        RECT 165.270 1.660 165.720 1.770 ;
        RECT 163.420 1.420 165.720 1.660 ;
        RECT 163.420 1.320 163.870 1.420 ;
        RECT 164.260 0.990 164.670 1.420 ;
        RECT 165.270 1.350 165.720 1.420 ;
        RECT 166.670 1.660 167.120 1.740 ;
        RECT 167.720 1.660 168.130 2.100 ;
        RECT 168.520 1.660 168.970 1.770 ;
        RECT 166.670 1.420 168.970 1.660 ;
        RECT 166.670 1.320 167.120 1.420 ;
        RECT 168.520 1.320 168.970 1.420 ;
        RECT 170.160 1.660 170.610 1.770 ;
        RECT 171.000 1.660 171.410 2.100 ;
        RECT 174.180 1.830 174.630 2.110 ;
        RECT 178.000 1.830 178.450 2.110 ;
        RECT 187.680 2.110 189.210 2.320 ;
        RECT 189.590 2.230 190.040 2.320 ;
        RECT 190.420 2.110 191.950 2.320 ;
        RECT 172.010 1.660 172.460 1.740 ;
        RECT 170.160 1.420 172.460 1.660 ;
        RECT 170.160 1.320 170.610 1.420 ;
        RECT 172.010 1.320 172.460 1.420 ;
        RECT 173.410 1.660 173.860 1.770 ;
        RECT 175.260 1.660 175.710 1.770 ;
        RECT 173.410 1.420 175.710 1.660 ;
        RECT 173.410 1.350 173.860 1.420 ;
        RECT 156.660 0.790 157.110 0.840 ;
        RECT 155.020 0.500 157.110 0.790 ;
        RECT 155.020 0.450 155.470 0.500 ;
        RECT 138.270 -0.130 138.720 -0.060 ;
        RECT 136.420 -0.370 138.720 -0.130 ;
        RECT 136.420 -0.480 136.870 -0.370 ;
        RECT 138.270 -0.480 138.720 -0.370 ;
        RECT 139.670 -0.130 140.120 -0.030 ;
        RECT 141.520 -0.130 141.970 -0.030 ;
        RECT 139.670 -0.370 141.970 -0.130 ;
        RECT 139.670 -0.450 140.120 -0.370 ;
        RECT 120.180 -1.030 121.710 -0.820 ;
        RECT 122.090 -1.030 122.540 -0.940 ;
        RECT 122.920 -1.030 124.450 -0.820 ;
        RECT 133.680 -0.820 134.130 -0.540 ;
        RECT 137.500 -0.820 137.950 -0.540 ;
        RECT 140.720 -0.810 141.130 -0.370 ;
        RECT 141.520 -0.480 141.970 -0.370 ;
        RECT 143.160 -0.130 143.610 -0.030 ;
        RECT 145.010 -0.130 145.460 -0.030 ;
        RECT 143.160 -0.370 145.460 -0.130 ;
        RECT 143.160 -0.480 143.610 -0.370 ;
        RECT 144.000 -0.810 144.410 -0.370 ;
        RECT 145.010 -0.450 145.460 -0.370 ;
        RECT 146.410 -0.130 146.860 -0.060 ;
        RECT 147.460 -0.130 147.870 0.300 ;
        RECT 148.260 -0.130 148.710 -0.030 ;
        RECT 146.410 -0.370 148.710 -0.130 ;
        RECT 146.410 -0.480 146.860 -0.370 ;
        RECT 148.260 -0.480 148.710 -0.370 ;
        RECT 149.920 -0.130 150.370 -0.030 ;
        RECT 150.760 -0.130 151.170 0.300 ;
        RECT 153.920 0.230 155.470 0.450 ;
        RECT 155.850 0.440 156.280 0.500 ;
        RECT 156.660 0.450 157.110 0.500 ;
        RECT 157.710 0.450 158.210 0.840 ;
        RECT 156.660 0.230 158.210 0.450 ;
        RECT 167.420 0.840 168.970 1.060 ;
        RECT 167.420 0.450 167.920 0.840 ;
        RECT 168.520 0.790 168.970 0.840 ;
        RECT 169.350 0.790 169.780 0.850 ;
        RECT 170.160 0.840 171.710 1.060 ;
        RECT 174.460 0.990 174.870 1.420 ;
        RECT 175.260 1.320 175.710 1.420 ;
        RECT 176.920 1.660 177.370 1.770 ;
        RECT 178.770 1.660 179.220 1.770 ;
        RECT 176.920 1.420 179.220 1.660 ;
        RECT 176.920 1.320 177.370 1.420 ;
        RECT 177.760 0.990 178.170 1.420 ;
        RECT 178.770 1.350 179.220 1.420 ;
        RECT 180.170 1.660 180.620 1.740 ;
        RECT 181.220 1.660 181.630 2.100 ;
        RECT 182.020 1.660 182.470 1.770 ;
        RECT 180.170 1.420 182.470 1.660 ;
        RECT 180.170 1.320 180.620 1.420 ;
        RECT 182.020 1.320 182.470 1.420 ;
        RECT 183.660 1.660 184.110 1.770 ;
        RECT 184.500 1.660 184.910 2.100 ;
        RECT 187.680 1.830 188.130 2.110 ;
        RECT 191.500 1.830 191.950 2.110 ;
        RECT 201.180 2.110 202.710 2.320 ;
        RECT 203.090 2.230 203.540 2.320 ;
        RECT 203.920 2.110 205.450 2.320 ;
        RECT 185.510 1.660 185.960 1.740 ;
        RECT 183.660 1.420 185.960 1.660 ;
        RECT 183.660 1.320 184.110 1.420 ;
        RECT 185.510 1.320 185.960 1.420 ;
        RECT 186.910 1.660 187.360 1.770 ;
        RECT 188.760 1.660 189.210 1.770 ;
        RECT 186.910 1.420 189.210 1.660 ;
        RECT 186.910 1.350 187.360 1.420 ;
        RECT 170.160 0.790 170.610 0.840 ;
        RECT 168.520 0.500 170.610 0.790 ;
        RECT 168.520 0.450 168.970 0.500 ;
        RECT 151.770 -0.130 152.220 -0.060 ;
        RECT 149.920 -0.370 152.220 -0.130 ;
        RECT 149.920 -0.480 150.370 -0.370 ;
        RECT 151.770 -0.480 152.220 -0.370 ;
        RECT 153.170 -0.130 153.620 -0.030 ;
        RECT 155.020 -0.130 155.470 -0.030 ;
        RECT 153.170 -0.370 155.470 -0.130 ;
        RECT 153.170 -0.450 153.620 -0.370 ;
        RECT 133.680 -1.030 135.210 -0.820 ;
        RECT 135.590 -1.030 136.040 -0.940 ;
        RECT 136.420 -1.030 137.950 -0.820 ;
        RECT 147.180 -0.820 147.630 -0.540 ;
        RECT 151.000 -0.820 151.450 -0.540 ;
        RECT 154.220 -0.810 154.630 -0.370 ;
        RECT 155.020 -0.480 155.470 -0.370 ;
        RECT 156.660 -0.130 157.110 -0.030 ;
        RECT 158.510 -0.130 158.960 -0.030 ;
        RECT 156.660 -0.370 158.960 -0.130 ;
        RECT 156.660 -0.480 157.110 -0.370 ;
        RECT 157.500 -0.810 157.910 -0.370 ;
        RECT 158.510 -0.450 158.960 -0.370 ;
        RECT 159.910 -0.130 160.360 -0.060 ;
        RECT 160.960 -0.130 161.370 0.300 ;
        RECT 161.760 -0.130 162.210 -0.030 ;
        RECT 159.910 -0.370 162.210 -0.130 ;
        RECT 159.910 -0.480 160.360 -0.370 ;
        RECT 161.760 -0.480 162.210 -0.370 ;
        RECT 163.420 -0.130 163.870 -0.030 ;
        RECT 164.260 -0.130 164.670 0.300 ;
        RECT 167.420 0.230 168.970 0.450 ;
        RECT 169.350 0.440 169.780 0.500 ;
        RECT 170.160 0.450 170.610 0.500 ;
        RECT 171.210 0.450 171.710 0.840 ;
        RECT 170.160 0.230 171.710 0.450 ;
        RECT 180.920 0.840 182.470 1.060 ;
        RECT 180.920 0.450 181.420 0.840 ;
        RECT 182.020 0.790 182.470 0.840 ;
        RECT 182.850 0.790 183.280 0.850 ;
        RECT 183.660 0.840 185.210 1.060 ;
        RECT 187.960 0.990 188.370 1.420 ;
        RECT 188.760 1.320 189.210 1.420 ;
        RECT 190.420 1.660 190.870 1.770 ;
        RECT 192.270 1.660 192.720 1.770 ;
        RECT 190.420 1.420 192.720 1.660 ;
        RECT 190.420 1.320 190.870 1.420 ;
        RECT 191.260 0.990 191.670 1.420 ;
        RECT 192.270 1.350 192.720 1.420 ;
        RECT 193.670 1.660 194.120 1.740 ;
        RECT 194.720 1.660 195.130 2.100 ;
        RECT 195.520 1.660 195.970 1.770 ;
        RECT 193.670 1.420 195.970 1.660 ;
        RECT 193.670 1.320 194.120 1.420 ;
        RECT 195.520 1.320 195.970 1.420 ;
        RECT 197.160 1.660 197.610 1.770 ;
        RECT 198.000 1.660 198.410 2.100 ;
        RECT 201.180 1.830 201.630 2.110 ;
        RECT 205.000 1.830 205.450 2.110 ;
        RECT 214.680 2.110 216.210 2.320 ;
        RECT 216.590 2.270 217.690 2.320 ;
        RECT 216.590 2.230 217.030 2.270 ;
        RECT 199.010 1.660 199.460 1.740 ;
        RECT 197.160 1.420 199.460 1.660 ;
        RECT 197.160 1.320 197.610 1.420 ;
        RECT 199.010 1.320 199.460 1.420 ;
        RECT 200.410 1.660 200.860 1.770 ;
        RECT 202.260 1.660 202.710 1.770 ;
        RECT 200.410 1.420 202.710 1.660 ;
        RECT 200.410 1.350 200.860 1.420 ;
        RECT 183.660 0.790 184.110 0.840 ;
        RECT 182.020 0.500 184.110 0.790 ;
        RECT 182.020 0.450 182.470 0.500 ;
        RECT 165.270 -0.130 165.720 -0.060 ;
        RECT 163.420 -0.370 165.720 -0.130 ;
        RECT 163.420 -0.480 163.870 -0.370 ;
        RECT 165.270 -0.480 165.720 -0.370 ;
        RECT 166.670 -0.130 167.120 -0.030 ;
        RECT 168.520 -0.130 168.970 -0.030 ;
        RECT 166.670 -0.370 168.970 -0.130 ;
        RECT 166.670 -0.450 167.120 -0.370 ;
        RECT 147.180 -1.030 148.710 -0.820 ;
        RECT 149.090 -1.030 149.540 -0.940 ;
        RECT 149.920 -1.030 151.450 -0.820 ;
        RECT 160.680 -0.820 161.130 -0.540 ;
        RECT 164.500 -0.820 164.950 -0.540 ;
        RECT 167.720 -0.810 168.130 -0.370 ;
        RECT 168.520 -0.480 168.970 -0.370 ;
        RECT 170.160 -0.130 170.610 -0.030 ;
        RECT 172.010 -0.130 172.460 -0.030 ;
        RECT 170.160 -0.370 172.460 -0.130 ;
        RECT 170.160 -0.480 170.610 -0.370 ;
        RECT 171.000 -0.810 171.410 -0.370 ;
        RECT 172.010 -0.450 172.460 -0.370 ;
        RECT 173.410 -0.130 173.860 -0.060 ;
        RECT 174.460 -0.130 174.870 0.300 ;
        RECT 175.260 -0.130 175.710 -0.030 ;
        RECT 173.410 -0.370 175.710 -0.130 ;
        RECT 173.410 -0.480 173.860 -0.370 ;
        RECT 175.260 -0.480 175.710 -0.370 ;
        RECT 176.920 -0.130 177.370 -0.030 ;
        RECT 177.760 -0.130 178.170 0.300 ;
        RECT 180.920 0.230 182.470 0.450 ;
        RECT 182.850 0.440 183.280 0.500 ;
        RECT 183.660 0.450 184.110 0.500 ;
        RECT 184.710 0.450 185.210 0.840 ;
        RECT 183.660 0.230 185.210 0.450 ;
        RECT 194.420 0.840 195.970 1.060 ;
        RECT 194.420 0.450 194.920 0.840 ;
        RECT 195.520 0.790 195.970 0.840 ;
        RECT 196.350 0.790 196.780 0.850 ;
        RECT 197.160 0.840 198.710 1.060 ;
        RECT 201.460 0.990 201.870 1.420 ;
        RECT 202.260 1.320 202.710 1.420 ;
        RECT 203.920 1.660 204.370 1.770 ;
        RECT 205.770 1.660 206.220 1.770 ;
        RECT 203.920 1.420 206.220 1.660 ;
        RECT 203.920 1.320 204.370 1.420 ;
        RECT 204.760 0.990 205.170 1.420 ;
        RECT 205.770 1.350 206.220 1.420 ;
        RECT 207.170 1.660 207.620 1.740 ;
        RECT 208.220 1.660 208.630 2.100 ;
        RECT 209.020 1.660 209.470 1.770 ;
        RECT 207.170 1.420 209.470 1.660 ;
        RECT 207.170 1.320 207.620 1.420 ;
        RECT 209.020 1.320 209.470 1.420 ;
        RECT 210.660 1.660 211.110 1.770 ;
        RECT 211.500 1.660 211.910 2.100 ;
        RECT 214.680 1.830 215.130 2.110 ;
        RECT 212.510 1.660 212.960 1.740 ;
        RECT 210.660 1.420 212.960 1.660 ;
        RECT 210.660 1.320 211.110 1.420 ;
        RECT 212.510 1.320 212.960 1.420 ;
        RECT 213.910 1.660 214.360 1.770 ;
        RECT 215.760 1.660 216.210 1.770 ;
        RECT 213.910 1.420 216.210 1.660 ;
        RECT 213.910 1.350 214.360 1.420 ;
        RECT 197.160 0.790 197.610 0.840 ;
        RECT 195.520 0.500 197.610 0.790 ;
        RECT 195.520 0.450 195.970 0.500 ;
        RECT 178.770 -0.130 179.220 -0.060 ;
        RECT 176.920 -0.370 179.220 -0.130 ;
        RECT 176.920 -0.480 177.370 -0.370 ;
        RECT 178.770 -0.480 179.220 -0.370 ;
        RECT 180.170 -0.130 180.620 -0.030 ;
        RECT 182.020 -0.130 182.470 -0.030 ;
        RECT 180.170 -0.370 182.470 -0.130 ;
        RECT 180.170 -0.450 180.620 -0.370 ;
        RECT 160.680 -1.030 162.210 -0.820 ;
        RECT 162.590 -1.030 163.040 -0.940 ;
        RECT 163.420 -1.030 164.950 -0.820 ;
        RECT 174.180 -0.820 174.630 -0.540 ;
        RECT 178.000 -0.820 178.450 -0.540 ;
        RECT 181.220 -0.810 181.630 -0.370 ;
        RECT 182.020 -0.480 182.470 -0.370 ;
        RECT 183.660 -0.130 184.110 -0.030 ;
        RECT 185.510 -0.130 185.960 -0.030 ;
        RECT 183.660 -0.370 185.960 -0.130 ;
        RECT 183.660 -0.480 184.110 -0.370 ;
        RECT 184.500 -0.810 184.910 -0.370 ;
        RECT 185.510 -0.450 185.960 -0.370 ;
        RECT 186.910 -0.130 187.360 -0.060 ;
        RECT 187.960 -0.130 188.370 0.300 ;
        RECT 188.760 -0.130 189.210 -0.030 ;
        RECT 186.910 -0.370 189.210 -0.130 ;
        RECT 186.910 -0.480 187.360 -0.370 ;
        RECT 188.760 -0.480 189.210 -0.370 ;
        RECT 190.420 -0.130 190.870 -0.030 ;
        RECT 191.260 -0.130 191.670 0.300 ;
        RECT 194.420 0.230 195.970 0.450 ;
        RECT 196.350 0.440 196.780 0.500 ;
        RECT 197.160 0.450 197.610 0.500 ;
        RECT 198.210 0.450 198.710 0.840 ;
        RECT 197.160 0.230 198.710 0.450 ;
        RECT 207.920 0.840 209.470 1.060 ;
        RECT 207.920 0.450 208.420 0.840 ;
        RECT 209.020 0.790 209.470 0.840 ;
        RECT 209.850 0.790 210.280 0.850 ;
        RECT 210.660 0.840 212.210 1.060 ;
        RECT 214.960 0.990 215.370 1.420 ;
        RECT 215.760 1.320 216.210 1.420 ;
        RECT 210.660 0.790 211.110 0.840 ;
        RECT 209.020 0.500 211.110 0.790 ;
        RECT 209.020 0.450 209.470 0.500 ;
        RECT 192.270 -0.130 192.720 -0.060 ;
        RECT 190.420 -0.370 192.720 -0.130 ;
        RECT 190.420 -0.480 190.870 -0.370 ;
        RECT 192.270 -0.480 192.720 -0.370 ;
        RECT 193.670 -0.130 194.120 -0.030 ;
        RECT 195.520 -0.130 195.970 -0.030 ;
        RECT 193.670 -0.370 195.970 -0.130 ;
        RECT 193.670 -0.450 194.120 -0.370 ;
        RECT 174.180 -1.030 175.710 -0.820 ;
        RECT 176.090 -1.030 176.540 -0.940 ;
        RECT 176.920 -1.030 178.450 -0.820 ;
        RECT 187.680 -0.820 188.130 -0.540 ;
        RECT 191.500 -0.820 191.950 -0.540 ;
        RECT 194.720 -0.810 195.130 -0.370 ;
        RECT 195.520 -0.480 195.970 -0.370 ;
        RECT 197.160 -0.130 197.610 -0.030 ;
        RECT 199.010 -0.130 199.460 -0.030 ;
        RECT 197.160 -0.370 199.460 -0.130 ;
        RECT 197.160 -0.480 197.610 -0.370 ;
        RECT 198.000 -0.810 198.410 -0.370 ;
        RECT 199.010 -0.450 199.460 -0.370 ;
        RECT 200.410 -0.130 200.860 -0.060 ;
        RECT 201.460 -0.130 201.870 0.300 ;
        RECT 202.260 -0.130 202.710 -0.030 ;
        RECT 200.410 -0.370 202.710 -0.130 ;
        RECT 200.410 -0.480 200.860 -0.370 ;
        RECT 202.260 -0.480 202.710 -0.370 ;
        RECT 203.920 -0.130 204.370 -0.030 ;
        RECT 204.760 -0.130 205.170 0.300 ;
        RECT 207.920 0.230 209.470 0.450 ;
        RECT 209.850 0.440 210.280 0.500 ;
        RECT 210.660 0.450 211.110 0.500 ;
        RECT 211.710 0.450 212.210 0.840 ;
        RECT 210.660 0.230 212.210 0.450 ;
        RECT 205.770 -0.130 206.220 -0.060 ;
        RECT 203.920 -0.370 206.220 -0.130 ;
        RECT 203.920 -0.480 204.370 -0.370 ;
        RECT 205.770 -0.480 206.220 -0.370 ;
        RECT 207.170 -0.130 207.620 -0.030 ;
        RECT 209.020 -0.130 209.470 -0.030 ;
        RECT 207.170 -0.370 209.470 -0.130 ;
        RECT 207.170 -0.450 207.620 -0.370 ;
        RECT 187.680 -1.030 189.210 -0.820 ;
        RECT 189.590 -1.030 190.040 -0.940 ;
        RECT 190.420 -1.030 191.950 -0.820 ;
        RECT 201.180 -0.820 201.630 -0.540 ;
        RECT 205.000 -0.820 205.450 -0.540 ;
        RECT 208.220 -0.810 208.630 -0.370 ;
        RECT 209.020 -0.480 209.470 -0.370 ;
        RECT 210.660 -0.130 211.110 -0.030 ;
        RECT 212.510 -0.130 212.960 -0.030 ;
        RECT 210.660 -0.370 212.960 -0.130 ;
        RECT 210.660 -0.480 211.110 -0.370 ;
        RECT 211.500 -0.810 211.910 -0.370 ;
        RECT 212.510 -0.450 212.960 -0.370 ;
        RECT 213.910 -0.130 214.360 -0.060 ;
        RECT 214.960 -0.130 215.370 0.300 ;
        RECT 215.760 -0.130 216.210 -0.030 ;
        RECT 213.910 -0.370 216.210 -0.130 ;
        RECT 213.910 -0.480 214.360 -0.370 ;
        RECT 215.760 -0.480 216.210 -0.370 ;
        RECT 201.180 -1.030 202.710 -0.820 ;
        RECT 203.090 -1.030 203.540 -0.940 ;
        RECT 203.920 -1.030 205.450 -0.820 ;
        RECT 214.680 -0.820 215.130 -0.540 ;
        RECT 214.680 -1.030 216.210 -0.820 ;
        RECT 216.590 -1.030 217.030 -0.940 ;
        RECT 13.260 -1.290 15.370 -1.030 ;
        RECT 26.760 -1.290 28.870 -1.030 ;
        RECT 40.260 -1.290 42.370 -1.030 ;
        RECT 53.760 -1.290 55.870 -1.030 ;
        RECT 67.260 -1.290 69.370 -1.030 ;
        RECT 80.760 -1.290 82.870 -1.030 ;
        RECT 94.260 -1.290 96.370 -1.030 ;
        RECT 107.760 -1.290 109.870 -1.030 ;
        RECT 121.260 -1.290 123.370 -1.030 ;
        RECT 134.760 -1.290 136.870 -1.030 ;
        RECT 148.260 -1.290 150.370 -1.030 ;
        RECT 161.760 -1.290 163.870 -1.030 ;
        RECT 175.260 -1.290 177.370 -1.030 ;
        RECT 188.760 -1.290 190.870 -1.030 ;
        RECT 202.260 -1.290 204.370 -1.030 ;
        RECT 215.760 -1.040 217.030 -1.030 ;
        RECT 215.760 -1.230 217.240 -1.040 ;
        RECT 215.760 -1.290 217.030 -1.230 ;
        RECT 12.180 -1.500 13.710 -1.290 ;
        RECT 14.090 -1.380 14.540 -1.290 ;
        RECT 14.920 -1.500 16.450 -1.290 ;
        RECT 1.420 -1.950 1.870 -1.840 ;
        RECT 3.270 -1.950 3.720 -1.840 ;
        RECT 1.420 -2.190 3.720 -1.950 ;
        RECT 1.420 -2.290 1.870 -2.190 ;
        RECT 2.260 -2.620 2.670 -2.190 ;
        RECT 3.270 -2.260 3.720 -2.190 ;
        RECT 4.670 -1.950 5.120 -1.870 ;
        RECT 5.720 -1.950 6.130 -1.510 ;
        RECT 6.520 -1.950 6.970 -1.840 ;
        RECT 4.670 -2.190 6.970 -1.950 ;
        RECT 4.670 -2.290 5.120 -2.190 ;
        RECT 6.520 -2.290 6.970 -2.190 ;
        RECT 8.160 -1.950 8.610 -1.840 ;
        RECT 9.000 -1.950 9.410 -1.510 ;
        RECT 12.180 -1.780 12.630 -1.500 ;
        RECT 16.000 -1.780 16.450 -1.500 ;
        RECT 25.680 -1.500 27.210 -1.290 ;
        RECT 27.590 -1.380 28.040 -1.290 ;
        RECT 28.420 -1.500 29.950 -1.290 ;
        RECT 10.010 -1.950 10.460 -1.870 ;
        RECT 8.160 -2.190 10.460 -1.950 ;
        RECT 8.160 -2.290 8.610 -2.190 ;
        RECT 10.010 -2.290 10.460 -2.190 ;
        RECT 11.410 -1.950 11.860 -1.840 ;
        RECT 13.260 -1.950 13.710 -1.840 ;
        RECT 11.410 -2.190 13.710 -1.950 ;
        RECT 11.410 -2.260 11.860 -2.190 ;
        RECT 5.420 -2.770 6.970 -2.550 ;
        RECT 5.420 -3.160 5.920 -2.770 ;
        RECT 6.520 -2.820 6.970 -2.770 ;
        RECT 7.350 -2.820 7.780 -2.760 ;
        RECT 8.160 -2.770 9.710 -2.550 ;
        RECT 12.460 -2.620 12.870 -2.190 ;
        RECT 13.260 -2.290 13.710 -2.190 ;
        RECT 14.920 -1.950 15.370 -1.840 ;
        RECT 16.770 -1.950 17.220 -1.840 ;
        RECT 14.920 -2.190 17.220 -1.950 ;
        RECT 14.920 -2.290 15.370 -2.190 ;
        RECT 15.760 -2.620 16.170 -2.190 ;
        RECT 16.770 -2.260 17.220 -2.190 ;
        RECT 18.170 -1.950 18.620 -1.870 ;
        RECT 19.220 -1.950 19.630 -1.510 ;
        RECT 20.020 -1.950 20.470 -1.840 ;
        RECT 18.170 -2.190 20.470 -1.950 ;
        RECT 18.170 -2.290 18.620 -2.190 ;
        RECT 20.020 -2.290 20.470 -2.190 ;
        RECT 21.660 -1.950 22.110 -1.840 ;
        RECT 22.500 -1.950 22.910 -1.510 ;
        RECT 25.680 -1.780 26.130 -1.500 ;
        RECT 29.500 -1.780 29.950 -1.500 ;
        RECT 39.180 -1.500 40.710 -1.290 ;
        RECT 41.090 -1.380 41.540 -1.290 ;
        RECT 41.920 -1.500 43.450 -1.290 ;
        RECT 23.510 -1.950 23.960 -1.870 ;
        RECT 21.660 -2.190 23.960 -1.950 ;
        RECT 21.660 -2.290 22.110 -2.190 ;
        RECT 23.510 -2.290 23.960 -2.190 ;
        RECT 24.910 -1.950 25.360 -1.840 ;
        RECT 26.760 -1.950 27.210 -1.840 ;
        RECT 24.910 -2.190 27.210 -1.950 ;
        RECT 24.910 -2.260 25.360 -2.190 ;
        RECT 8.160 -2.820 8.610 -2.770 ;
        RECT 6.520 -3.110 8.610 -2.820 ;
        RECT 6.520 -3.160 6.970 -3.110 ;
        RECT 1.420 -3.740 1.870 -3.640 ;
        RECT 2.260 -3.740 2.670 -3.310 ;
        RECT 5.420 -3.380 6.970 -3.160 ;
        RECT 7.350 -3.170 7.780 -3.110 ;
        RECT 8.160 -3.160 8.610 -3.110 ;
        RECT 9.210 -3.160 9.710 -2.770 ;
        RECT 8.160 -3.380 9.710 -3.160 ;
        RECT 18.920 -2.770 20.470 -2.550 ;
        RECT 18.920 -3.160 19.420 -2.770 ;
        RECT 20.020 -2.820 20.470 -2.770 ;
        RECT 20.850 -2.820 21.280 -2.760 ;
        RECT 21.660 -2.770 23.210 -2.550 ;
        RECT 25.960 -2.620 26.370 -2.190 ;
        RECT 26.760 -2.290 27.210 -2.190 ;
        RECT 28.420 -1.950 28.870 -1.840 ;
        RECT 30.270 -1.950 30.720 -1.840 ;
        RECT 28.420 -2.190 30.720 -1.950 ;
        RECT 28.420 -2.290 28.870 -2.190 ;
        RECT 29.260 -2.620 29.670 -2.190 ;
        RECT 30.270 -2.260 30.720 -2.190 ;
        RECT 31.670 -1.950 32.120 -1.870 ;
        RECT 32.720 -1.950 33.130 -1.510 ;
        RECT 33.520 -1.950 33.970 -1.840 ;
        RECT 31.670 -2.190 33.970 -1.950 ;
        RECT 31.670 -2.290 32.120 -2.190 ;
        RECT 33.520 -2.290 33.970 -2.190 ;
        RECT 35.160 -1.950 35.610 -1.840 ;
        RECT 36.000 -1.950 36.410 -1.510 ;
        RECT 39.180 -1.780 39.630 -1.500 ;
        RECT 43.000 -1.780 43.450 -1.500 ;
        RECT 52.680 -1.500 54.210 -1.290 ;
        RECT 54.590 -1.380 55.040 -1.290 ;
        RECT 55.420 -1.500 56.950 -1.290 ;
        RECT 37.010 -1.950 37.460 -1.870 ;
        RECT 35.160 -2.190 37.460 -1.950 ;
        RECT 35.160 -2.290 35.610 -2.190 ;
        RECT 37.010 -2.290 37.460 -2.190 ;
        RECT 38.410 -1.950 38.860 -1.840 ;
        RECT 40.260 -1.950 40.710 -1.840 ;
        RECT 38.410 -2.190 40.710 -1.950 ;
        RECT 38.410 -2.260 38.860 -2.190 ;
        RECT 21.660 -2.820 22.110 -2.770 ;
        RECT 20.020 -3.110 22.110 -2.820 ;
        RECT 20.020 -3.160 20.470 -3.110 ;
        RECT 3.270 -3.740 3.720 -3.670 ;
        RECT 1.420 -3.980 3.720 -3.740 ;
        RECT 1.420 -4.090 1.870 -3.980 ;
        RECT 3.270 -4.090 3.720 -3.980 ;
        RECT 4.670 -3.740 5.120 -3.640 ;
        RECT 6.520 -3.740 6.970 -3.640 ;
        RECT 4.670 -3.980 6.970 -3.740 ;
        RECT 4.670 -4.060 5.120 -3.980 ;
        RECT 5.720 -4.420 6.130 -3.980 ;
        RECT 6.520 -4.090 6.970 -3.980 ;
        RECT 8.160 -3.740 8.610 -3.640 ;
        RECT 10.010 -3.740 10.460 -3.640 ;
        RECT 8.160 -3.980 10.460 -3.740 ;
        RECT 8.160 -4.090 8.610 -3.980 ;
        RECT 9.000 -4.420 9.410 -3.980 ;
        RECT 10.010 -4.060 10.460 -3.980 ;
        RECT 11.410 -3.740 11.860 -3.670 ;
        RECT 12.460 -3.740 12.870 -3.310 ;
        RECT 13.260 -3.740 13.710 -3.640 ;
        RECT 11.410 -3.980 13.710 -3.740 ;
        RECT 11.410 -4.090 11.860 -3.980 ;
        RECT 13.260 -4.090 13.710 -3.980 ;
        RECT 14.920 -3.740 15.370 -3.640 ;
        RECT 15.760 -3.740 16.170 -3.310 ;
        RECT 18.920 -3.380 20.470 -3.160 ;
        RECT 20.850 -3.170 21.280 -3.110 ;
        RECT 21.660 -3.160 22.110 -3.110 ;
        RECT 22.710 -3.160 23.210 -2.770 ;
        RECT 21.660 -3.380 23.210 -3.160 ;
        RECT 32.420 -2.770 33.970 -2.550 ;
        RECT 32.420 -3.160 32.920 -2.770 ;
        RECT 33.520 -2.820 33.970 -2.770 ;
        RECT 34.350 -2.820 34.780 -2.760 ;
        RECT 35.160 -2.770 36.710 -2.550 ;
        RECT 39.460 -2.620 39.870 -2.190 ;
        RECT 40.260 -2.290 40.710 -2.190 ;
        RECT 41.920 -1.950 42.370 -1.840 ;
        RECT 43.770 -1.950 44.220 -1.840 ;
        RECT 41.920 -2.190 44.220 -1.950 ;
        RECT 41.920 -2.290 42.370 -2.190 ;
        RECT 42.760 -2.620 43.170 -2.190 ;
        RECT 43.770 -2.260 44.220 -2.190 ;
        RECT 45.170 -1.950 45.620 -1.870 ;
        RECT 46.220 -1.950 46.630 -1.510 ;
        RECT 47.020 -1.950 47.470 -1.840 ;
        RECT 45.170 -2.190 47.470 -1.950 ;
        RECT 45.170 -2.290 45.620 -2.190 ;
        RECT 47.020 -2.290 47.470 -2.190 ;
        RECT 48.660 -1.950 49.110 -1.840 ;
        RECT 49.500 -1.950 49.910 -1.510 ;
        RECT 52.680 -1.780 53.130 -1.500 ;
        RECT 56.500 -1.780 56.950 -1.500 ;
        RECT 66.180 -1.500 67.710 -1.290 ;
        RECT 68.090 -1.380 68.540 -1.290 ;
        RECT 68.920 -1.500 70.450 -1.290 ;
        RECT 50.510 -1.950 50.960 -1.870 ;
        RECT 48.660 -2.190 50.960 -1.950 ;
        RECT 48.660 -2.290 49.110 -2.190 ;
        RECT 50.510 -2.290 50.960 -2.190 ;
        RECT 51.910 -1.950 52.360 -1.840 ;
        RECT 53.760 -1.950 54.210 -1.840 ;
        RECT 51.910 -2.190 54.210 -1.950 ;
        RECT 51.910 -2.260 52.360 -2.190 ;
        RECT 35.160 -2.820 35.610 -2.770 ;
        RECT 33.520 -3.110 35.610 -2.820 ;
        RECT 33.520 -3.160 33.970 -3.110 ;
        RECT 16.770 -3.740 17.220 -3.670 ;
        RECT 14.920 -3.980 17.220 -3.740 ;
        RECT 14.920 -4.090 15.370 -3.980 ;
        RECT 16.770 -4.090 17.220 -3.980 ;
        RECT 18.170 -3.740 18.620 -3.640 ;
        RECT 20.020 -3.740 20.470 -3.640 ;
        RECT 18.170 -3.980 20.470 -3.740 ;
        RECT 18.170 -4.060 18.620 -3.980 ;
        RECT 12.180 -4.430 12.630 -4.150 ;
        RECT 16.000 -4.430 16.450 -4.150 ;
        RECT 19.220 -4.420 19.630 -3.980 ;
        RECT 20.020 -4.090 20.470 -3.980 ;
        RECT 21.660 -3.740 22.110 -3.640 ;
        RECT 23.510 -3.740 23.960 -3.640 ;
        RECT 21.660 -3.980 23.960 -3.740 ;
        RECT 21.660 -4.090 22.110 -3.980 ;
        RECT 22.500 -4.420 22.910 -3.980 ;
        RECT 23.510 -4.060 23.960 -3.980 ;
        RECT 24.910 -3.740 25.360 -3.670 ;
        RECT 25.960 -3.740 26.370 -3.310 ;
        RECT 26.760 -3.740 27.210 -3.640 ;
        RECT 24.910 -3.980 27.210 -3.740 ;
        RECT 24.910 -4.090 25.360 -3.980 ;
        RECT 26.760 -4.090 27.210 -3.980 ;
        RECT 28.420 -3.740 28.870 -3.640 ;
        RECT 29.260 -3.740 29.670 -3.310 ;
        RECT 32.420 -3.380 33.970 -3.160 ;
        RECT 34.350 -3.170 34.780 -3.110 ;
        RECT 35.160 -3.160 35.610 -3.110 ;
        RECT 36.210 -3.160 36.710 -2.770 ;
        RECT 35.160 -3.380 36.710 -3.160 ;
        RECT 45.920 -2.770 47.470 -2.550 ;
        RECT 45.920 -3.160 46.420 -2.770 ;
        RECT 47.020 -2.820 47.470 -2.770 ;
        RECT 47.850 -2.820 48.280 -2.760 ;
        RECT 48.660 -2.770 50.210 -2.550 ;
        RECT 52.960 -2.620 53.370 -2.190 ;
        RECT 53.760 -2.290 54.210 -2.190 ;
        RECT 55.420 -1.950 55.870 -1.840 ;
        RECT 57.270 -1.950 57.720 -1.840 ;
        RECT 55.420 -2.190 57.720 -1.950 ;
        RECT 55.420 -2.290 55.870 -2.190 ;
        RECT 56.260 -2.620 56.670 -2.190 ;
        RECT 57.270 -2.260 57.720 -2.190 ;
        RECT 58.670 -1.950 59.120 -1.870 ;
        RECT 59.720 -1.950 60.130 -1.510 ;
        RECT 60.520 -1.950 60.970 -1.840 ;
        RECT 58.670 -2.190 60.970 -1.950 ;
        RECT 58.670 -2.290 59.120 -2.190 ;
        RECT 60.520 -2.290 60.970 -2.190 ;
        RECT 62.160 -1.950 62.610 -1.840 ;
        RECT 63.000 -1.950 63.410 -1.510 ;
        RECT 66.180 -1.780 66.630 -1.500 ;
        RECT 70.000 -1.780 70.450 -1.500 ;
        RECT 79.680 -1.500 81.210 -1.290 ;
        RECT 81.590 -1.380 82.040 -1.290 ;
        RECT 82.420 -1.500 83.950 -1.290 ;
        RECT 64.010 -1.950 64.460 -1.870 ;
        RECT 62.160 -2.190 64.460 -1.950 ;
        RECT 62.160 -2.290 62.610 -2.190 ;
        RECT 64.010 -2.290 64.460 -2.190 ;
        RECT 65.410 -1.950 65.860 -1.840 ;
        RECT 67.260 -1.950 67.710 -1.840 ;
        RECT 65.410 -2.190 67.710 -1.950 ;
        RECT 65.410 -2.260 65.860 -2.190 ;
        RECT 48.660 -2.820 49.110 -2.770 ;
        RECT 47.020 -3.110 49.110 -2.820 ;
        RECT 47.020 -3.160 47.470 -3.110 ;
        RECT 30.270 -3.740 30.720 -3.670 ;
        RECT 28.420 -3.980 30.720 -3.740 ;
        RECT 28.420 -4.090 28.870 -3.980 ;
        RECT 30.270 -4.090 30.720 -3.980 ;
        RECT 31.670 -3.740 32.120 -3.640 ;
        RECT 33.520 -3.740 33.970 -3.640 ;
        RECT 31.670 -3.980 33.970 -3.740 ;
        RECT 31.670 -4.060 32.120 -3.980 ;
        RECT 12.180 -4.640 13.710 -4.430 ;
        RECT 14.090 -4.640 14.540 -4.550 ;
        RECT 14.920 -4.640 16.450 -4.430 ;
        RECT 25.680 -4.430 26.130 -4.150 ;
        RECT 29.500 -4.430 29.950 -4.150 ;
        RECT 32.720 -4.420 33.130 -3.980 ;
        RECT 33.520 -4.090 33.970 -3.980 ;
        RECT 35.160 -3.740 35.610 -3.640 ;
        RECT 37.010 -3.740 37.460 -3.640 ;
        RECT 35.160 -3.980 37.460 -3.740 ;
        RECT 35.160 -4.090 35.610 -3.980 ;
        RECT 36.000 -4.420 36.410 -3.980 ;
        RECT 37.010 -4.060 37.460 -3.980 ;
        RECT 38.410 -3.740 38.860 -3.670 ;
        RECT 39.460 -3.740 39.870 -3.310 ;
        RECT 40.260 -3.740 40.710 -3.640 ;
        RECT 38.410 -3.980 40.710 -3.740 ;
        RECT 38.410 -4.090 38.860 -3.980 ;
        RECT 40.260 -4.090 40.710 -3.980 ;
        RECT 41.920 -3.740 42.370 -3.640 ;
        RECT 42.760 -3.740 43.170 -3.310 ;
        RECT 45.920 -3.380 47.470 -3.160 ;
        RECT 47.850 -3.170 48.280 -3.110 ;
        RECT 48.660 -3.160 49.110 -3.110 ;
        RECT 49.710 -3.160 50.210 -2.770 ;
        RECT 48.660 -3.380 50.210 -3.160 ;
        RECT 59.420 -2.770 60.970 -2.550 ;
        RECT 59.420 -3.160 59.920 -2.770 ;
        RECT 60.520 -2.820 60.970 -2.770 ;
        RECT 61.350 -2.820 61.780 -2.760 ;
        RECT 62.160 -2.770 63.710 -2.550 ;
        RECT 66.460 -2.620 66.870 -2.190 ;
        RECT 67.260 -2.290 67.710 -2.190 ;
        RECT 68.920 -1.950 69.370 -1.840 ;
        RECT 70.770 -1.950 71.220 -1.840 ;
        RECT 68.920 -2.190 71.220 -1.950 ;
        RECT 68.920 -2.290 69.370 -2.190 ;
        RECT 69.760 -2.620 70.170 -2.190 ;
        RECT 70.770 -2.260 71.220 -2.190 ;
        RECT 72.170 -1.950 72.620 -1.870 ;
        RECT 73.220 -1.950 73.630 -1.510 ;
        RECT 74.020 -1.950 74.470 -1.840 ;
        RECT 72.170 -2.190 74.470 -1.950 ;
        RECT 72.170 -2.290 72.620 -2.190 ;
        RECT 74.020 -2.290 74.470 -2.190 ;
        RECT 75.660 -1.950 76.110 -1.840 ;
        RECT 76.500 -1.950 76.910 -1.510 ;
        RECT 79.680 -1.780 80.130 -1.500 ;
        RECT 83.500 -1.780 83.950 -1.500 ;
        RECT 93.180 -1.500 94.710 -1.290 ;
        RECT 95.090 -1.380 95.540 -1.290 ;
        RECT 95.920 -1.500 97.450 -1.290 ;
        RECT 77.510 -1.950 77.960 -1.870 ;
        RECT 75.660 -2.190 77.960 -1.950 ;
        RECT 75.660 -2.290 76.110 -2.190 ;
        RECT 77.510 -2.290 77.960 -2.190 ;
        RECT 78.910 -1.950 79.360 -1.840 ;
        RECT 80.760 -1.950 81.210 -1.840 ;
        RECT 78.910 -2.190 81.210 -1.950 ;
        RECT 78.910 -2.260 79.360 -2.190 ;
        RECT 62.160 -2.820 62.610 -2.770 ;
        RECT 60.520 -3.110 62.610 -2.820 ;
        RECT 60.520 -3.160 60.970 -3.110 ;
        RECT 43.770 -3.740 44.220 -3.670 ;
        RECT 41.920 -3.980 44.220 -3.740 ;
        RECT 41.920 -4.090 42.370 -3.980 ;
        RECT 43.770 -4.090 44.220 -3.980 ;
        RECT 45.170 -3.740 45.620 -3.640 ;
        RECT 47.020 -3.740 47.470 -3.640 ;
        RECT 45.170 -3.980 47.470 -3.740 ;
        RECT 45.170 -4.060 45.620 -3.980 ;
        RECT 25.680 -4.640 27.210 -4.430 ;
        RECT 27.590 -4.640 28.040 -4.550 ;
        RECT 28.420 -4.640 29.950 -4.430 ;
        RECT 39.180 -4.430 39.630 -4.150 ;
        RECT 43.000 -4.430 43.450 -4.150 ;
        RECT 46.220 -4.420 46.630 -3.980 ;
        RECT 47.020 -4.090 47.470 -3.980 ;
        RECT 48.660 -3.740 49.110 -3.640 ;
        RECT 50.510 -3.740 50.960 -3.640 ;
        RECT 48.660 -3.980 50.960 -3.740 ;
        RECT 48.660 -4.090 49.110 -3.980 ;
        RECT 49.500 -4.420 49.910 -3.980 ;
        RECT 50.510 -4.060 50.960 -3.980 ;
        RECT 51.910 -3.740 52.360 -3.670 ;
        RECT 52.960 -3.740 53.370 -3.310 ;
        RECT 53.760 -3.740 54.210 -3.640 ;
        RECT 51.910 -3.980 54.210 -3.740 ;
        RECT 51.910 -4.090 52.360 -3.980 ;
        RECT 53.760 -4.090 54.210 -3.980 ;
        RECT 55.420 -3.740 55.870 -3.640 ;
        RECT 56.260 -3.740 56.670 -3.310 ;
        RECT 59.420 -3.380 60.970 -3.160 ;
        RECT 61.350 -3.170 61.780 -3.110 ;
        RECT 62.160 -3.160 62.610 -3.110 ;
        RECT 63.210 -3.160 63.710 -2.770 ;
        RECT 62.160 -3.380 63.710 -3.160 ;
        RECT 72.920 -2.770 74.470 -2.550 ;
        RECT 72.920 -3.160 73.420 -2.770 ;
        RECT 74.020 -2.820 74.470 -2.770 ;
        RECT 74.850 -2.820 75.280 -2.760 ;
        RECT 75.660 -2.770 77.210 -2.550 ;
        RECT 79.960 -2.620 80.370 -2.190 ;
        RECT 80.760 -2.290 81.210 -2.190 ;
        RECT 82.420 -1.950 82.870 -1.840 ;
        RECT 84.270 -1.950 84.720 -1.840 ;
        RECT 82.420 -2.190 84.720 -1.950 ;
        RECT 82.420 -2.290 82.870 -2.190 ;
        RECT 83.260 -2.620 83.670 -2.190 ;
        RECT 84.270 -2.260 84.720 -2.190 ;
        RECT 85.670 -1.950 86.120 -1.870 ;
        RECT 86.720 -1.950 87.130 -1.510 ;
        RECT 87.520 -1.950 87.970 -1.840 ;
        RECT 85.670 -2.190 87.970 -1.950 ;
        RECT 85.670 -2.290 86.120 -2.190 ;
        RECT 87.520 -2.290 87.970 -2.190 ;
        RECT 89.160 -1.950 89.610 -1.840 ;
        RECT 90.000 -1.950 90.410 -1.510 ;
        RECT 93.180 -1.780 93.630 -1.500 ;
        RECT 97.000 -1.780 97.450 -1.500 ;
        RECT 106.680 -1.500 108.210 -1.290 ;
        RECT 108.590 -1.380 109.040 -1.290 ;
        RECT 109.420 -1.500 110.950 -1.290 ;
        RECT 91.010 -1.950 91.460 -1.870 ;
        RECT 89.160 -2.190 91.460 -1.950 ;
        RECT 89.160 -2.290 89.610 -2.190 ;
        RECT 91.010 -2.290 91.460 -2.190 ;
        RECT 92.410 -1.950 92.860 -1.840 ;
        RECT 94.260 -1.950 94.710 -1.840 ;
        RECT 92.410 -2.190 94.710 -1.950 ;
        RECT 92.410 -2.260 92.860 -2.190 ;
        RECT 75.660 -2.820 76.110 -2.770 ;
        RECT 74.020 -3.110 76.110 -2.820 ;
        RECT 74.020 -3.160 74.470 -3.110 ;
        RECT 57.270 -3.740 57.720 -3.670 ;
        RECT 55.420 -3.980 57.720 -3.740 ;
        RECT 55.420 -4.090 55.870 -3.980 ;
        RECT 57.270 -4.090 57.720 -3.980 ;
        RECT 58.670 -3.740 59.120 -3.640 ;
        RECT 60.520 -3.740 60.970 -3.640 ;
        RECT 58.670 -3.980 60.970 -3.740 ;
        RECT 58.670 -4.060 59.120 -3.980 ;
        RECT 39.180 -4.640 40.710 -4.430 ;
        RECT 41.090 -4.640 41.540 -4.550 ;
        RECT 41.920 -4.640 43.450 -4.430 ;
        RECT 52.680 -4.430 53.130 -4.150 ;
        RECT 56.500 -4.430 56.950 -4.150 ;
        RECT 59.720 -4.420 60.130 -3.980 ;
        RECT 60.520 -4.090 60.970 -3.980 ;
        RECT 62.160 -3.740 62.610 -3.640 ;
        RECT 64.010 -3.740 64.460 -3.640 ;
        RECT 62.160 -3.980 64.460 -3.740 ;
        RECT 62.160 -4.090 62.610 -3.980 ;
        RECT 63.000 -4.420 63.410 -3.980 ;
        RECT 64.010 -4.060 64.460 -3.980 ;
        RECT 65.410 -3.740 65.860 -3.670 ;
        RECT 66.460 -3.740 66.870 -3.310 ;
        RECT 67.260 -3.740 67.710 -3.640 ;
        RECT 65.410 -3.980 67.710 -3.740 ;
        RECT 65.410 -4.090 65.860 -3.980 ;
        RECT 67.260 -4.090 67.710 -3.980 ;
        RECT 68.920 -3.740 69.370 -3.640 ;
        RECT 69.760 -3.740 70.170 -3.310 ;
        RECT 72.920 -3.380 74.470 -3.160 ;
        RECT 74.850 -3.170 75.280 -3.110 ;
        RECT 75.660 -3.160 76.110 -3.110 ;
        RECT 76.710 -3.160 77.210 -2.770 ;
        RECT 75.660 -3.380 77.210 -3.160 ;
        RECT 86.420 -2.770 87.970 -2.550 ;
        RECT 86.420 -3.160 86.920 -2.770 ;
        RECT 87.520 -2.820 87.970 -2.770 ;
        RECT 88.350 -2.820 88.780 -2.760 ;
        RECT 89.160 -2.770 90.710 -2.550 ;
        RECT 93.460 -2.620 93.870 -2.190 ;
        RECT 94.260 -2.290 94.710 -2.190 ;
        RECT 95.920 -1.950 96.370 -1.840 ;
        RECT 97.770 -1.950 98.220 -1.840 ;
        RECT 95.920 -2.190 98.220 -1.950 ;
        RECT 95.920 -2.290 96.370 -2.190 ;
        RECT 96.760 -2.620 97.170 -2.190 ;
        RECT 97.770 -2.260 98.220 -2.190 ;
        RECT 99.170 -1.950 99.620 -1.870 ;
        RECT 100.220 -1.950 100.630 -1.510 ;
        RECT 101.020 -1.950 101.470 -1.840 ;
        RECT 99.170 -2.190 101.470 -1.950 ;
        RECT 99.170 -2.290 99.620 -2.190 ;
        RECT 101.020 -2.290 101.470 -2.190 ;
        RECT 102.660 -1.950 103.110 -1.840 ;
        RECT 103.500 -1.950 103.910 -1.510 ;
        RECT 106.680 -1.780 107.130 -1.500 ;
        RECT 110.500 -1.780 110.950 -1.500 ;
        RECT 120.180 -1.500 121.710 -1.290 ;
        RECT 122.090 -1.380 122.540 -1.290 ;
        RECT 122.920 -1.500 124.450 -1.290 ;
        RECT 104.510 -1.950 104.960 -1.870 ;
        RECT 102.660 -2.190 104.960 -1.950 ;
        RECT 102.660 -2.290 103.110 -2.190 ;
        RECT 104.510 -2.290 104.960 -2.190 ;
        RECT 105.910 -1.950 106.360 -1.840 ;
        RECT 107.760 -1.950 108.210 -1.840 ;
        RECT 105.910 -2.190 108.210 -1.950 ;
        RECT 105.910 -2.260 106.360 -2.190 ;
        RECT 89.160 -2.820 89.610 -2.770 ;
        RECT 87.520 -3.110 89.610 -2.820 ;
        RECT 87.520 -3.160 87.970 -3.110 ;
        RECT 70.770 -3.740 71.220 -3.670 ;
        RECT 68.920 -3.980 71.220 -3.740 ;
        RECT 68.920 -4.090 69.370 -3.980 ;
        RECT 70.770 -4.090 71.220 -3.980 ;
        RECT 72.170 -3.740 72.620 -3.640 ;
        RECT 74.020 -3.740 74.470 -3.640 ;
        RECT 72.170 -3.980 74.470 -3.740 ;
        RECT 72.170 -4.060 72.620 -3.980 ;
        RECT 52.680 -4.640 54.210 -4.430 ;
        RECT 54.590 -4.640 55.040 -4.550 ;
        RECT 55.420 -4.640 56.950 -4.430 ;
        RECT 66.180 -4.430 66.630 -4.150 ;
        RECT 70.000 -4.430 70.450 -4.150 ;
        RECT 73.220 -4.420 73.630 -3.980 ;
        RECT 74.020 -4.090 74.470 -3.980 ;
        RECT 75.660 -3.740 76.110 -3.640 ;
        RECT 77.510 -3.740 77.960 -3.640 ;
        RECT 75.660 -3.980 77.960 -3.740 ;
        RECT 75.660 -4.090 76.110 -3.980 ;
        RECT 76.500 -4.420 76.910 -3.980 ;
        RECT 77.510 -4.060 77.960 -3.980 ;
        RECT 78.910 -3.740 79.360 -3.670 ;
        RECT 79.960 -3.740 80.370 -3.310 ;
        RECT 80.760 -3.740 81.210 -3.640 ;
        RECT 78.910 -3.980 81.210 -3.740 ;
        RECT 78.910 -4.090 79.360 -3.980 ;
        RECT 80.760 -4.090 81.210 -3.980 ;
        RECT 82.420 -3.740 82.870 -3.640 ;
        RECT 83.260 -3.740 83.670 -3.310 ;
        RECT 86.420 -3.380 87.970 -3.160 ;
        RECT 88.350 -3.170 88.780 -3.110 ;
        RECT 89.160 -3.160 89.610 -3.110 ;
        RECT 90.210 -3.160 90.710 -2.770 ;
        RECT 89.160 -3.380 90.710 -3.160 ;
        RECT 99.920 -2.770 101.470 -2.550 ;
        RECT 99.920 -3.160 100.420 -2.770 ;
        RECT 101.020 -2.820 101.470 -2.770 ;
        RECT 101.850 -2.820 102.280 -2.760 ;
        RECT 102.660 -2.770 104.210 -2.550 ;
        RECT 106.960 -2.620 107.370 -2.190 ;
        RECT 107.760 -2.290 108.210 -2.190 ;
        RECT 109.420 -1.950 109.870 -1.840 ;
        RECT 111.270 -1.950 111.720 -1.840 ;
        RECT 109.420 -2.190 111.720 -1.950 ;
        RECT 109.420 -2.290 109.870 -2.190 ;
        RECT 110.260 -2.620 110.670 -2.190 ;
        RECT 111.270 -2.260 111.720 -2.190 ;
        RECT 112.670 -1.950 113.120 -1.870 ;
        RECT 113.720 -1.950 114.130 -1.510 ;
        RECT 114.520 -1.950 114.970 -1.840 ;
        RECT 112.670 -2.190 114.970 -1.950 ;
        RECT 112.670 -2.290 113.120 -2.190 ;
        RECT 114.520 -2.290 114.970 -2.190 ;
        RECT 116.160 -1.950 116.610 -1.840 ;
        RECT 117.000 -1.950 117.410 -1.510 ;
        RECT 120.180 -1.780 120.630 -1.500 ;
        RECT 124.000 -1.780 124.450 -1.500 ;
        RECT 133.680 -1.500 135.210 -1.290 ;
        RECT 135.590 -1.380 136.040 -1.290 ;
        RECT 136.420 -1.500 137.950 -1.290 ;
        RECT 118.010 -1.950 118.460 -1.870 ;
        RECT 116.160 -2.190 118.460 -1.950 ;
        RECT 116.160 -2.290 116.610 -2.190 ;
        RECT 118.010 -2.290 118.460 -2.190 ;
        RECT 119.410 -1.950 119.860 -1.840 ;
        RECT 121.260 -1.950 121.710 -1.840 ;
        RECT 119.410 -2.190 121.710 -1.950 ;
        RECT 119.410 -2.260 119.860 -2.190 ;
        RECT 102.660 -2.820 103.110 -2.770 ;
        RECT 101.020 -3.110 103.110 -2.820 ;
        RECT 101.020 -3.160 101.470 -3.110 ;
        RECT 84.270 -3.740 84.720 -3.670 ;
        RECT 82.420 -3.980 84.720 -3.740 ;
        RECT 82.420 -4.090 82.870 -3.980 ;
        RECT 84.270 -4.090 84.720 -3.980 ;
        RECT 85.670 -3.740 86.120 -3.640 ;
        RECT 87.520 -3.740 87.970 -3.640 ;
        RECT 85.670 -3.980 87.970 -3.740 ;
        RECT 85.670 -4.060 86.120 -3.980 ;
        RECT 66.180 -4.640 67.710 -4.430 ;
        RECT 68.090 -4.640 68.540 -4.550 ;
        RECT 68.920 -4.640 70.450 -4.430 ;
        RECT 79.680 -4.430 80.130 -4.150 ;
        RECT 83.500 -4.430 83.950 -4.150 ;
        RECT 86.720 -4.420 87.130 -3.980 ;
        RECT 87.520 -4.090 87.970 -3.980 ;
        RECT 89.160 -3.740 89.610 -3.640 ;
        RECT 91.010 -3.740 91.460 -3.640 ;
        RECT 89.160 -3.980 91.460 -3.740 ;
        RECT 89.160 -4.090 89.610 -3.980 ;
        RECT 90.000 -4.420 90.410 -3.980 ;
        RECT 91.010 -4.060 91.460 -3.980 ;
        RECT 92.410 -3.740 92.860 -3.670 ;
        RECT 93.460 -3.740 93.870 -3.310 ;
        RECT 94.260 -3.740 94.710 -3.640 ;
        RECT 92.410 -3.980 94.710 -3.740 ;
        RECT 92.410 -4.090 92.860 -3.980 ;
        RECT 94.260 -4.090 94.710 -3.980 ;
        RECT 95.920 -3.740 96.370 -3.640 ;
        RECT 96.760 -3.740 97.170 -3.310 ;
        RECT 99.920 -3.380 101.470 -3.160 ;
        RECT 101.850 -3.170 102.280 -3.110 ;
        RECT 102.660 -3.160 103.110 -3.110 ;
        RECT 103.710 -3.160 104.210 -2.770 ;
        RECT 102.660 -3.380 104.210 -3.160 ;
        RECT 113.420 -2.770 114.970 -2.550 ;
        RECT 113.420 -3.160 113.920 -2.770 ;
        RECT 114.520 -2.820 114.970 -2.770 ;
        RECT 115.350 -2.820 115.780 -2.760 ;
        RECT 116.160 -2.770 117.710 -2.550 ;
        RECT 120.460 -2.620 120.870 -2.190 ;
        RECT 121.260 -2.290 121.710 -2.190 ;
        RECT 122.920 -1.950 123.370 -1.840 ;
        RECT 124.770 -1.950 125.220 -1.840 ;
        RECT 122.920 -2.190 125.220 -1.950 ;
        RECT 122.920 -2.290 123.370 -2.190 ;
        RECT 123.760 -2.620 124.170 -2.190 ;
        RECT 124.770 -2.260 125.220 -2.190 ;
        RECT 126.170 -1.950 126.620 -1.870 ;
        RECT 127.220 -1.950 127.630 -1.510 ;
        RECT 128.020 -1.950 128.470 -1.840 ;
        RECT 126.170 -2.190 128.470 -1.950 ;
        RECT 126.170 -2.290 126.620 -2.190 ;
        RECT 128.020 -2.290 128.470 -2.190 ;
        RECT 129.660 -1.950 130.110 -1.840 ;
        RECT 130.500 -1.950 130.910 -1.510 ;
        RECT 133.680 -1.780 134.130 -1.500 ;
        RECT 137.500 -1.780 137.950 -1.500 ;
        RECT 147.180 -1.500 148.710 -1.290 ;
        RECT 149.090 -1.380 149.540 -1.290 ;
        RECT 149.920 -1.500 151.450 -1.290 ;
        RECT 131.510 -1.950 131.960 -1.870 ;
        RECT 129.660 -2.190 131.960 -1.950 ;
        RECT 129.660 -2.290 130.110 -2.190 ;
        RECT 131.510 -2.290 131.960 -2.190 ;
        RECT 132.910 -1.950 133.360 -1.840 ;
        RECT 134.760 -1.950 135.210 -1.840 ;
        RECT 132.910 -2.190 135.210 -1.950 ;
        RECT 132.910 -2.260 133.360 -2.190 ;
        RECT 116.160 -2.820 116.610 -2.770 ;
        RECT 114.520 -3.110 116.610 -2.820 ;
        RECT 114.520 -3.160 114.970 -3.110 ;
        RECT 97.770 -3.740 98.220 -3.670 ;
        RECT 95.920 -3.980 98.220 -3.740 ;
        RECT 95.920 -4.090 96.370 -3.980 ;
        RECT 97.770 -4.090 98.220 -3.980 ;
        RECT 99.170 -3.740 99.620 -3.640 ;
        RECT 101.020 -3.740 101.470 -3.640 ;
        RECT 99.170 -3.980 101.470 -3.740 ;
        RECT 99.170 -4.060 99.620 -3.980 ;
        RECT 79.680 -4.640 81.210 -4.430 ;
        RECT 81.590 -4.640 82.040 -4.550 ;
        RECT 82.420 -4.640 83.950 -4.430 ;
        RECT 93.180 -4.430 93.630 -4.150 ;
        RECT 97.000 -4.430 97.450 -4.150 ;
        RECT 100.220 -4.420 100.630 -3.980 ;
        RECT 101.020 -4.090 101.470 -3.980 ;
        RECT 102.660 -3.740 103.110 -3.640 ;
        RECT 104.510 -3.740 104.960 -3.640 ;
        RECT 102.660 -3.980 104.960 -3.740 ;
        RECT 102.660 -4.090 103.110 -3.980 ;
        RECT 103.500 -4.420 103.910 -3.980 ;
        RECT 104.510 -4.060 104.960 -3.980 ;
        RECT 105.910 -3.740 106.360 -3.670 ;
        RECT 106.960 -3.740 107.370 -3.310 ;
        RECT 107.760 -3.740 108.210 -3.640 ;
        RECT 105.910 -3.980 108.210 -3.740 ;
        RECT 105.910 -4.090 106.360 -3.980 ;
        RECT 107.760 -4.090 108.210 -3.980 ;
        RECT 109.420 -3.740 109.870 -3.640 ;
        RECT 110.260 -3.740 110.670 -3.310 ;
        RECT 113.420 -3.380 114.970 -3.160 ;
        RECT 115.350 -3.170 115.780 -3.110 ;
        RECT 116.160 -3.160 116.610 -3.110 ;
        RECT 117.210 -3.160 117.710 -2.770 ;
        RECT 116.160 -3.380 117.710 -3.160 ;
        RECT 126.920 -2.770 128.470 -2.550 ;
        RECT 126.920 -3.160 127.420 -2.770 ;
        RECT 128.020 -2.820 128.470 -2.770 ;
        RECT 128.850 -2.820 129.280 -2.760 ;
        RECT 129.660 -2.770 131.210 -2.550 ;
        RECT 133.960 -2.620 134.370 -2.190 ;
        RECT 134.760 -2.290 135.210 -2.190 ;
        RECT 136.420 -1.950 136.870 -1.840 ;
        RECT 138.270 -1.950 138.720 -1.840 ;
        RECT 136.420 -2.190 138.720 -1.950 ;
        RECT 136.420 -2.290 136.870 -2.190 ;
        RECT 137.260 -2.620 137.670 -2.190 ;
        RECT 138.270 -2.260 138.720 -2.190 ;
        RECT 139.670 -1.950 140.120 -1.870 ;
        RECT 140.720 -1.950 141.130 -1.510 ;
        RECT 141.520 -1.950 141.970 -1.840 ;
        RECT 139.670 -2.190 141.970 -1.950 ;
        RECT 139.670 -2.290 140.120 -2.190 ;
        RECT 141.520 -2.290 141.970 -2.190 ;
        RECT 143.160 -1.950 143.610 -1.840 ;
        RECT 144.000 -1.950 144.410 -1.510 ;
        RECT 147.180 -1.780 147.630 -1.500 ;
        RECT 151.000 -1.780 151.450 -1.500 ;
        RECT 160.680 -1.500 162.210 -1.290 ;
        RECT 162.590 -1.380 163.040 -1.290 ;
        RECT 163.420 -1.500 164.950 -1.290 ;
        RECT 145.010 -1.950 145.460 -1.870 ;
        RECT 143.160 -2.190 145.460 -1.950 ;
        RECT 143.160 -2.290 143.610 -2.190 ;
        RECT 145.010 -2.290 145.460 -2.190 ;
        RECT 146.410 -1.950 146.860 -1.840 ;
        RECT 148.260 -1.950 148.710 -1.840 ;
        RECT 146.410 -2.190 148.710 -1.950 ;
        RECT 146.410 -2.260 146.860 -2.190 ;
        RECT 129.660 -2.820 130.110 -2.770 ;
        RECT 128.020 -3.110 130.110 -2.820 ;
        RECT 128.020 -3.160 128.470 -3.110 ;
        RECT 111.270 -3.740 111.720 -3.670 ;
        RECT 109.420 -3.980 111.720 -3.740 ;
        RECT 109.420 -4.090 109.870 -3.980 ;
        RECT 111.270 -4.090 111.720 -3.980 ;
        RECT 112.670 -3.740 113.120 -3.640 ;
        RECT 114.520 -3.740 114.970 -3.640 ;
        RECT 112.670 -3.980 114.970 -3.740 ;
        RECT 112.670 -4.060 113.120 -3.980 ;
        RECT 93.180 -4.640 94.710 -4.430 ;
        RECT 95.090 -4.640 95.540 -4.550 ;
        RECT 95.920 -4.640 97.450 -4.430 ;
        RECT 106.680 -4.430 107.130 -4.150 ;
        RECT 110.500 -4.430 110.950 -4.150 ;
        RECT 113.720 -4.420 114.130 -3.980 ;
        RECT 114.520 -4.090 114.970 -3.980 ;
        RECT 116.160 -3.740 116.610 -3.640 ;
        RECT 118.010 -3.740 118.460 -3.640 ;
        RECT 116.160 -3.980 118.460 -3.740 ;
        RECT 116.160 -4.090 116.610 -3.980 ;
        RECT 117.000 -4.420 117.410 -3.980 ;
        RECT 118.010 -4.060 118.460 -3.980 ;
        RECT 119.410 -3.740 119.860 -3.670 ;
        RECT 120.460 -3.740 120.870 -3.310 ;
        RECT 121.260 -3.740 121.710 -3.640 ;
        RECT 119.410 -3.980 121.710 -3.740 ;
        RECT 119.410 -4.090 119.860 -3.980 ;
        RECT 121.260 -4.090 121.710 -3.980 ;
        RECT 122.920 -3.740 123.370 -3.640 ;
        RECT 123.760 -3.740 124.170 -3.310 ;
        RECT 126.920 -3.380 128.470 -3.160 ;
        RECT 128.850 -3.170 129.280 -3.110 ;
        RECT 129.660 -3.160 130.110 -3.110 ;
        RECT 130.710 -3.160 131.210 -2.770 ;
        RECT 129.660 -3.380 131.210 -3.160 ;
        RECT 140.420 -2.770 141.970 -2.550 ;
        RECT 140.420 -3.160 140.920 -2.770 ;
        RECT 141.520 -2.820 141.970 -2.770 ;
        RECT 142.350 -2.820 142.780 -2.760 ;
        RECT 143.160 -2.770 144.710 -2.550 ;
        RECT 147.460 -2.620 147.870 -2.190 ;
        RECT 148.260 -2.290 148.710 -2.190 ;
        RECT 149.920 -1.950 150.370 -1.840 ;
        RECT 151.770 -1.950 152.220 -1.840 ;
        RECT 149.920 -2.190 152.220 -1.950 ;
        RECT 149.920 -2.290 150.370 -2.190 ;
        RECT 150.760 -2.620 151.170 -2.190 ;
        RECT 151.770 -2.260 152.220 -2.190 ;
        RECT 153.170 -1.950 153.620 -1.870 ;
        RECT 154.220 -1.950 154.630 -1.510 ;
        RECT 155.020 -1.950 155.470 -1.840 ;
        RECT 153.170 -2.190 155.470 -1.950 ;
        RECT 153.170 -2.290 153.620 -2.190 ;
        RECT 155.020 -2.290 155.470 -2.190 ;
        RECT 156.660 -1.950 157.110 -1.840 ;
        RECT 157.500 -1.950 157.910 -1.510 ;
        RECT 160.680 -1.780 161.130 -1.500 ;
        RECT 164.500 -1.780 164.950 -1.500 ;
        RECT 174.180 -1.500 175.710 -1.290 ;
        RECT 176.090 -1.380 176.540 -1.290 ;
        RECT 176.920 -1.500 178.450 -1.290 ;
        RECT 158.510 -1.950 158.960 -1.870 ;
        RECT 156.660 -2.190 158.960 -1.950 ;
        RECT 156.660 -2.290 157.110 -2.190 ;
        RECT 158.510 -2.290 158.960 -2.190 ;
        RECT 159.910 -1.950 160.360 -1.840 ;
        RECT 161.760 -1.950 162.210 -1.840 ;
        RECT 159.910 -2.190 162.210 -1.950 ;
        RECT 159.910 -2.260 160.360 -2.190 ;
        RECT 143.160 -2.820 143.610 -2.770 ;
        RECT 141.520 -3.110 143.610 -2.820 ;
        RECT 141.520 -3.160 141.970 -3.110 ;
        RECT 124.770 -3.740 125.220 -3.670 ;
        RECT 122.920 -3.980 125.220 -3.740 ;
        RECT 122.920 -4.090 123.370 -3.980 ;
        RECT 124.770 -4.090 125.220 -3.980 ;
        RECT 126.170 -3.740 126.620 -3.640 ;
        RECT 128.020 -3.740 128.470 -3.640 ;
        RECT 126.170 -3.980 128.470 -3.740 ;
        RECT 126.170 -4.060 126.620 -3.980 ;
        RECT 106.680 -4.640 108.210 -4.430 ;
        RECT 108.590 -4.640 109.040 -4.550 ;
        RECT 109.420 -4.640 110.950 -4.430 ;
        RECT 120.180 -4.430 120.630 -4.150 ;
        RECT 124.000 -4.430 124.450 -4.150 ;
        RECT 127.220 -4.420 127.630 -3.980 ;
        RECT 128.020 -4.090 128.470 -3.980 ;
        RECT 129.660 -3.740 130.110 -3.640 ;
        RECT 131.510 -3.740 131.960 -3.640 ;
        RECT 129.660 -3.980 131.960 -3.740 ;
        RECT 129.660 -4.090 130.110 -3.980 ;
        RECT 130.500 -4.420 130.910 -3.980 ;
        RECT 131.510 -4.060 131.960 -3.980 ;
        RECT 132.910 -3.740 133.360 -3.670 ;
        RECT 133.960 -3.740 134.370 -3.310 ;
        RECT 134.760 -3.740 135.210 -3.640 ;
        RECT 132.910 -3.980 135.210 -3.740 ;
        RECT 132.910 -4.090 133.360 -3.980 ;
        RECT 134.760 -4.090 135.210 -3.980 ;
        RECT 136.420 -3.740 136.870 -3.640 ;
        RECT 137.260 -3.740 137.670 -3.310 ;
        RECT 140.420 -3.380 141.970 -3.160 ;
        RECT 142.350 -3.170 142.780 -3.110 ;
        RECT 143.160 -3.160 143.610 -3.110 ;
        RECT 144.210 -3.160 144.710 -2.770 ;
        RECT 143.160 -3.380 144.710 -3.160 ;
        RECT 153.920 -2.770 155.470 -2.550 ;
        RECT 153.920 -3.160 154.420 -2.770 ;
        RECT 155.020 -2.820 155.470 -2.770 ;
        RECT 155.850 -2.820 156.280 -2.760 ;
        RECT 156.660 -2.770 158.210 -2.550 ;
        RECT 160.960 -2.620 161.370 -2.190 ;
        RECT 161.760 -2.290 162.210 -2.190 ;
        RECT 163.420 -1.950 163.870 -1.840 ;
        RECT 165.270 -1.950 165.720 -1.840 ;
        RECT 163.420 -2.190 165.720 -1.950 ;
        RECT 163.420 -2.290 163.870 -2.190 ;
        RECT 164.260 -2.620 164.670 -2.190 ;
        RECT 165.270 -2.260 165.720 -2.190 ;
        RECT 166.670 -1.950 167.120 -1.870 ;
        RECT 167.720 -1.950 168.130 -1.510 ;
        RECT 168.520 -1.950 168.970 -1.840 ;
        RECT 166.670 -2.190 168.970 -1.950 ;
        RECT 166.670 -2.290 167.120 -2.190 ;
        RECT 168.520 -2.290 168.970 -2.190 ;
        RECT 170.160 -1.950 170.610 -1.840 ;
        RECT 171.000 -1.950 171.410 -1.510 ;
        RECT 174.180 -1.780 174.630 -1.500 ;
        RECT 178.000 -1.780 178.450 -1.500 ;
        RECT 187.680 -1.500 189.210 -1.290 ;
        RECT 189.590 -1.380 190.040 -1.290 ;
        RECT 190.420 -1.500 191.950 -1.290 ;
        RECT 172.010 -1.950 172.460 -1.870 ;
        RECT 170.160 -2.190 172.460 -1.950 ;
        RECT 170.160 -2.290 170.610 -2.190 ;
        RECT 172.010 -2.290 172.460 -2.190 ;
        RECT 173.410 -1.950 173.860 -1.840 ;
        RECT 175.260 -1.950 175.710 -1.840 ;
        RECT 173.410 -2.190 175.710 -1.950 ;
        RECT 173.410 -2.260 173.860 -2.190 ;
        RECT 156.660 -2.820 157.110 -2.770 ;
        RECT 155.020 -3.110 157.110 -2.820 ;
        RECT 155.020 -3.160 155.470 -3.110 ;
        RECT 138.270 -3.740 138.720 -3.670 ;
        RECT 136.420 -3.980 138.720 -3.740 ;
        RECT 136.420 -4.090 136.870 -3.980 ;
        RECT 138.270 -4.090 138.720 -3.980 ;
        RECT 139.670 -3.740 140.120 -3.640 ;
        RECT 141.520 -3.740 141.970 -3.640 ;
        RECT 139.670 -3.980 141.970 -3.740 ;
        RECT 139.670 -4.060 140.120 -3.980 ;
        RECT 120.180 -4.640 121.710 -4.430 ;
        RECT 122.090 -4.640 122.540 -4.550 ;
        RECT 122.920 -4.640 124.450 -4.430 ;
        RECT 133.680 -4.430 134.130 -4.150 ;
        RECT 137.500 -4.430 137.950 -4.150 ;
        RECT 140.720 -4.420 141.130 -3.980 ;
        RECT 141.520 -4.090 141.970 -3.980 ;
        RECT 143.160 -3.740 143.610 -3.640 ;
        RECT 145.010 -3.740 145.460 -3.640 ;
        RECT 143.160 -3.980 145.460 -3.740 ;
        RECT 143.160 -4.090 143.610 -3.980 ;
        RECT 144.000 -4.420 144.410 -3.980 ;
        RECT 145.010 -4.060 145.460 -3.980 ;
        RECT 146.410 -3.740 146.860 -3.670 ;
        RECT 147.460 -3.740 147.870 -3.310 ;
        RECT 148.260 -3.740 148.710 -3.640 ;
        RECT 146.410 -3.980 148.710 -3.740 ;
        RECT 146.410 -4.090 146.860 -3.980 ;
        RECT 148.260 -4.090 148.710 -3.980 ;
        RECT 149.920 -3.740 150.370 -3.640 ;
        RECT 150.760 -3.740 151.170 -3.310 ;
        RECT 153.920 -3.380 155.470 -3.160 ;
        RECT 155.850 -3.170 156.280 -3.110 ;
        RECT 156.660 -3.160 157.110 -3.110 ;
        RECT 157.710 -3.160 158.210 -2.770 ;
        RECT 156.660 -3.380 158.210 -3.160 ;
        RECT 167.420 -2.770 168.970 -2.550 ;
        RECT 167.420 -3.160 167.920 -2.770 ;
        RECT 168.520 -2.820 168.970 -2.770 ;
        RECT 169.350 -2.820 169.780 -2.760 ;
        RECT 170.160 -2.770 171.710 -2.550 ;
        RECT 174.460 -2.620 174.870 -2.190 ;
        RECT 175.260 -2.290 175.710 -2.190 ;
        RECT 176.920 -1.950 177.370 -1.840 ;
        RECT 178.770 -1.950 179.220 -1.840 ;
        RECT 176.920 -2.190 179.220 -1.950 ;
        RECT 176.920 -2.290 177.370 -2.190 ;
        RECT 177.760 -2.620 178.170 -2.190 ;
        RECT 178.770 -2.260 179.220 -2.190 ;
        RECT 180.170 -1.950 180.620 -1.870 ;
        RECT 181.220 -1.950 181.630 -1.510 ;
        RECT 182.020 -1.950 182.470 -1.840 ;
        RECT 180.170 -2.190 182.470 -1.950 ;
        RECT 180.170 -2.290 180.620 -2.190 ;
        RECT 182.020 -2.290 182.470 -2.190 ;
        RECT 183.660 -1.950 184.110 -1.840 ;
        RECT 184.500 -1.950 184.910 -1.510 ;
        RECT 187.680 -1.780 188.130 -1.500 ;
        RECT 191.500 -1.780 191.950 -1.500 ;
        RECT 201.180 -1.500 202.710 -1.290 ;
        RECT 203.090 -1.380 203.540 -1.290 ;
        RECT 203.920 -1.500 205.450 -1.290 ;
        RECT 185.510 -1.950 185.960 -1.870 ;
        RECT 183.660 -2.190 185.960 -1.950 ;
        RECT 183.660 -2.290 184.110 -2.190 ;
        RECT 185.510 -2.290 185.960 -2.190 ;
        RECT 186.910 -1.950 187.360 -1.840 ;
        RECT 188.760 -1.950 189.210 -1.840 ;
        RECT 186.910 -2.190 189.210 -1.950 ;
        RECT 186.910 -2.260 187.360 -2.190 ;
        RECT 170.160 -2.820 170.610 -2.770 ;
        RECT 168.520 -3.110 170.610 -2.820 ;
        RECT 168.520 -3.160 168.970 -3.110 ;
        RECT 151.770 -3.740 152.220 -3.670 ;
        RECT 149.920 -3.980 152.220 -3.740 ;
        RECT 149.920 -4.090 150.370 -3.980 ;
        RECT 151.770 -4.090 152.220 -3.980 ;
        RECT 153.170 -3.740 153.620 -3.640 ;
        RECT 155.020 -3.740 155.470 -3.640 ;
        RECT 153.170 -3.980 155.470 -3.740 ;
        RECT 153.170 -4.060 153.620 -3.980 ;
        RECT 133.680 -4.640 135.210 -4.430 ;
        RECT 135.590 -4.640 136.040 -4.550 ;
        RECT 136.420 -4.640 137.950 -4.430 ;
        RECT 147.180 -4.430 147.630 -4.150 ;
        RECT 151.000 -4.430 151.450 -4.150 ;
        RECT 154.220 -4.420 154.630 -3.980 ;
        RECT 155.020 -4.090 155.470 -3.980 ;
        RECT 156.660 -3.740 157.110 -3.640 ;
        RECT 158.510 -3.740 158.960 -3.640 ;
        RECT 156.660 -3.980 158.960 -3.740 ;
        RECT 156.660 -4.090 157.110 -3.980 ;
        RECT 157.500 -4.420 157.910 -3.980 ;
        RECT 158.510 -4.060 158.960 -3.980 ;
        RECT 159.910 -3.740 160.360 -3.670 ;
        RECT 160.960 -3.740 161.370 -3.310 ;
        RECT 161.760 -3.740 162.210 -3.640 ;
        RECT 159.910 -3.980 162.210 -3.740 ;
        RECT 159.910 -4.090 160.360 -3.980 ;
        RECT 161.760 -4.090 162.210 -3.980 ;
        RECT 163.420 -3.740 163.870 -3.640 ;
        RECT 164.260 -3.740 164.670 -3.310 ;
        RECT 167.420 -3.380 168.970 -3.160 ;
        RECT 169.350 -3.170 169.780 -3.110 ;
        RECT 170.160 -3.160 170.610 -3.110 ;
        RECT 171.210 -3.160 171.710 -2.770 ;
        RECT 170.160 -3.380 171.710 -3.160 ;
        RECT 180.920 -2.770 182.470 -2.550 ;
        RECT 180.920 -3.160 181.420 -2.770 ;
        RECT 182.020 -2.820 182.470 -2.770 ;
        RECT 182.850 -2.820 183.280 -2.760 ;
        RECT 183.660 -2.770 185.210 -2.550 ;
        RECT 187.960 -2.620 188.370 -2.190 ;
        RECT 188.760 -2.290 189.210 -2.190 ;
        RECT 190.420 -1.950 190.870 -1.840 ;
        RECT 192.270 -1.950 192.720 -1.840 ;
        RECT 190.420 -2.190 192.720 -1.950 ;
        RECT 190.420 -2.290 190.870 -2.190 ;
        RECT 191.260 -2.620 191.670 -2.190 ;
        RECT 192.270 -2.260 192.720 -2.190 ;
        RECT 193.670 -1.950 194.120 -1.870 ;
        RECT 194.720 -1.950 195.130 -1.510 ;
        RECT 195.520 -1.950 195.970 -1.840 ;
        RECT 193.670 -2.190 195.970 -1.950 ;
        RECT 193.670 -2.290 194.120 -2.190 ;
        RECT 195.520 -2.290 195.970 -2.190 ;
        RECT 197.160 -1.950 197.610 -1.840 ;
        RECT 198.000 -1.950 198.410 -1.510 ;
        RECT 201.180 -1.780 201.630 -1.500 ;
        RECT 205.000 -1.780 205.450 -1.500 ;
        RECT 214.680 -1.500 216.210 -1.290 ;
        RECT 216.590 -1.380 217.030 -1.290 ;
        RECT 199.010 -1.950 199.460 -1.870 ;
        RECT 197.160 -2.190 199.460 -1.950 ;
        RECT 197.160 -2.290 197.610 -2.190 ;
        RECT 199.010 -2.290 199.460 -2.190 ;
        RECT 200.410 -1.950 200.860 -1.840 ;
        RECT 202.260 -1.950 202.710 -1.840 ;
        RECT 200.410 -2.190 202.710 -1.950 ;
        RECT 200.410 -2.260 200.860 -2.190 ;
        RECT 183.660 -2.820 184.110 -2.770 ;
        RECT 182.020 -3.110 184.110 -2.820 ;
        RECT 182.020 -3.160 182.470 -3.110 ;
        RECT 165.270 -3.740 165.720 -3.670 ;
        RECT 163.420 -3.980 165.720 -3.740 ;
        RECT 163.420 -4.090 163.870 -3.980 ;
        RECT 165.270 -4.090 165.720 -3.980 ;
        RECT 166.670 -3.740 167.120 -3.640 ;
        RECT 168.520 -3.740 168.970 -3.640 ;
        RECT 166.670 -3.980 168.970 -3.740 ;
        RECT 166.670 -4.060 167.120 -3.980 ;
        RECT 147.180 -4.640 148.710 -4.430 ;
        RECT 149.090 -4.640 149.540 -4.550 ;
        RECT 149.920 -4.640 151.450 -4.430 ;
        RECT 160.680 -4.430 161.130 -4.150 ;
        RECT 164.500 -4.430 164.950 -4.150 ;
        RECT 167.720 -4.420 168.130 -3.980 ;
        RECT 168.520 -4.090 168.970 -3.980 ;
        RECT 170.160 -3.740 170.610 -3.640 ;
        RECT 172.010 -3.740 172.460 -3.640 ;
        RECT 170.160 -3.980 172.460 -3.740 ;
        RECT 170.160 -4.090 170.610 -3.980 ;
        RECT 171.000 -4.420 171.410 -3.980 ;
        RECT 172.010 -4.060 172.460 -3.980 ;
        RECT 173.410 -3.740 173.860 -3.670 ;
        RECT 174.460 -3.740 174.870 -3.310 ;
        RECT 175.260 -3.740 175.710 -3.640 ;
        RECT 173.410 -3.980 175.710 -3.740 ;
        RECT 173.410 -4.090 173.860 -3.980 ;
        RECT 175.260 -4.090 175.710 -3.980 ;
        RECT 176.920 -3.740 177.370 -3.640 ;
        RECT 177.760 -3.740 178.170 -3.310 ;
        RECT 180.920 -3.380 182.470 -3.160 ;
        RECT 182.850 -3.170 183.280 -3.110 ;
        RECT 183.660 -3.160 184.110 -3.110 ;
        RECT 184.710 -3.160 185.210 -2.770 ;
        RECT 183.660 -3.380 185.210 -3.160 ;
        RECT 194.420 -2.770 195.970 -2.550 ;
        RECT 194.420 -3.160 194.920 -2.770 ;
        RECT 195.520 -2.820 195.970 -2.770 ;
        RECT 196.350 -2.820 196.780 -2.760 ;
        RECT 197.160 -2.770 198.710 -2.550 ;
        RECT 201.460 -2.620 201.870 -2.190 ;
        RECT 202.260 -2.290 202.710 -2.190 ;
        RECT 203.920 -1.950 204.370 -1.840 ;
        RECT 205.770 -1.950 206.220 -1.840 ;
        RECT 203.920 -2.190 206.220 -1.950 ;
        RECT 203.920 -2.290 204.370 -2.190 ;
        RECT 204.760 -2.620 205.170 -2.190 ;
        RECT 205.770 -2.260 206.220 -2.190 ;
        RECT 207.170 -1.950 207.620 -1.870 ;
        RECT 208.220 -1.950 208.630 -1.510 ;
        RECT 209.020 -1.950 209.470 -1.840 ;
        RECT 207.170 -2.190 209.470 -1.950 ;
        RECT 207.170 -2.290 207.620 -2.190 ;
        RECT 209.020 -2.290 209.470 -2.190 ;
        RECT 210.660 -1.950 211.110 -1.840 ;
        RECT 211.500 -1.950 211.910 -1.510 ;
        RECT 214.680 -1.780 215.130 -1.500 ;
        RECT 212.510 -1.950 212.960 -1.870 ;
        RECT 210.660 -2.190 212.960 -1.950 ;
        RECT 210.660 -2.290 211.110 -2.190 ;
        RECT 212.510 -2.290 212.960 -2.190 ;
        RECT 213.910 -1.950 214.360 -1.840 ;
        RECT 215.760 -1.950 216.210 -1.840 ;
        RECT 213.910 -2.190 216.210 -1.950 ;
        RECT 213.910 -2.260 214.360 -2.190 ;
        RECT 197.160 -2.820 197.610 -2.770 ;
        RECT 195.520 -3.110 197.610 -2.820 ;
        RECT 195.520 -3.160 195.970 -3.110 ;
        RECT 178.770 -3.740 179.220 -3.670 ;
        RECT 176.920 -3.980 179.220 -3.740 ;
        RECT 176.920 -4.090 177.370 -3.980 ;
        RECT 178.770 -4.090 179.220 -3.980 ;
        RECT 180.170 -3.740 180.620 -3.640 ;
        RECT 182.020 -3.740 182.470 -3.640 ;
        RECT 180.170 -3.980 182.470 -3.740 ;
        RECT 180.170 -4.060 180.620 -3.980 ;
        RECT 160.680 -4.640 162.210 -4.430 ;
        RECT 162.590 -4.640 163.040 -4.550 ;
        RECT 163.420 -4.640 164.950 -4.430 ;
        RECT 174.180 -4.430 174.630 -4.150 ;
        RECT 178.000 -4.430 178.450 -4.150 ;
        RECT 181.220 -4.420 181.630 -3.980 ;
        RECT 182.020 -4.090 182.470 -3.980 ;
        RECT 183.660 -3.740 184.110 -3.640 ;
        RECT 185.510 -3.740 185.960 -3.640 ;
        RECT 183.660 -3.980 185.960 -3.740 ;
        RECT 183.660 -4.090 184.110 -3.980 ;
        RECT 184.500 -4.420 184.910 -3.980 ;
        RECT 185.510 -4.060 185.960 -3.980 ;
        RECT 186.910 -3.740 187.360 -3.670 ;
        RECT 187.960 -3.740 188.370 -3.310 ;
        RECT 188.760 -3.740 189.210 -3.640 ;
        RECT 186.910 -3.980 189.210 -3.740 ;
        RECT 186.910 -4.090 187.360 -3.980 ;
        RECT 188.760 -4.090 189.210 -3.980 ;
        RECT 190.420 -3.740 190.870 -3.640 ;
        RECT 191.260 -3.740 191.670 -3.310 ;
        RECT 194.420 -3.380 195.970 -3.160 ;
        RECT 196.350 -3.170 196.780 -3.110 ;
        RECT 197.160 -3.160 197.610 -3.110 ;
        RECT 198.210 -3.160 198.710 -2.770 ;
        RECT 197.160 -3.380 198.710 -3.160 ;
        RECT 207.920 -2.770 209.470 -2.550 ;
        RECT 207.920 -3.160 208.420 -2.770 ;
        RECT 209.020 -2.820 209.470 -2.770 ;
        RECT 209.850 -2.820 210.280 -2.760 ;
        RECT 210.660 -2.770 212.210 -2.550 ;
        RECT 214.960 -2.620 215.370 -2.190 ;
        RECT 215.760 -2.290 216.210 -2.190 ;
        RECT 210.660 -2.820 211.110 -2.770 ;
        RECT 209.020 -3.110 211.110 -2.820 ;
        RECT 209.020 -3.160 209.470 -3.110 ;
        RECT 192.270 -3.740 192.720 -3.670 ;
        RECT 190.420 -3.980 192.720 -3.740 ;
        RECT 190.420 -4.090 190.870 -3.980 ;
        RECT 192.270 -4.090 192.720 -3.980 ;
        RECT 193.670 -3.740 194.120 -3.640 ;
        RECT 195.520 -3.740 195.970 -3.640 ;
        RECT 193.670 -3.980 195.970 -3.740 ;
        RECT 193.670 -4.060 194.120 -3.980 ;
        RECT 174.180 -4.640 175.710 -4.430 ;
        RECT 176.090 -4.640 176.540 -4.550 ;
        RECT 176.920 -4.640 178.450 -4.430 ;
        RECT 187.680 -4.430 188.130 -4.150 ;
        RECT 191.500 -4.430 191.950 -4.150 ;
        RECT 194.720 -4.420 195.130 -3.980 ;
        RECT 195.520 -4.090 195.970 -3.980 ;
        RECT 197.160 -3.740 197.610 -3.640 ;
        RECT 199.010 -3.740 199.460 -3.640 ;
        RECT 197.160 -3.980 199.460 -3.740 ;
        RECT 197.160 -4.090 197.610 -3.980 ;
        RECT 198.000 -4.420 198.410 -3.980 ;
        RECT 199.010 -4.060 199.460 -3.980 ;
        RECT 200.410 -3.740 200.860 -3.670 ;
        RECT 201.460 -3.740 201.870 -3.310 ;
        RECT 202.260 -3.740 202.710 -3.640 ;
        RECT 200.410 -3.980 202.710 -3.740 ;
        RECT 200.410 -4.090 200.860 -3.980 ;
        RECT 202.260 -4.090 202.710 -3.980 ;
        RECT 203.920 -3.740 204.370 -3.640 ;
        RECT 204.760 -3.740 205.170 -3.310 ;
        RECT 207.920 -3.380 209.470 -3.160 ;
        RECT 209.850 -3.170 210.280 -3.110 ;
        RECT 210.660 -3.160 211.110 -3.110 ;
        RECT 211.710 -3.160 212.210 -2.770 ;
        RECT 210.660 -3.380 212.210 -3.160 ;
        RECT 205.770 -3.740 206.220 -3.670 ;
        RECT 203.920 -3.980 206.220 -3.740 ;
        RECT 203.920 -4.090 204.370 -3.980 ;
        RECT 205.770 -4.090 206.220 -3.980 ;
        RECT 207.170 -3.740 207.620 -3.640 ;
        RECT 209.020 -3.740 209.470 -3.640 ;
        RECT 207.170 -3.980 209.470 -3.740 ;
        RECT 207.170 -4.060 207.620 -3.980 ;
        RECT 187.680 -4.640 189.210 -4.430 ;
        RECT 189.590 -4.640 190.040 -4.550 ;
        RECT 190.420 -4.640 191.950 -4.430 ;
        RECT 201.180 -4.430 201.630 -4.150 ;
        RECT 205.000 -4.430 205.450 -4.150 ;
        RECT 208.220 -4.420 208.630 -3.980 ;
        RECT 209.020 -4.090 209.470 -3.980 ;
        RECT 210.660 -3.740 211.110 -3.640 ;
        RECT 212.510 -3.740 212.960 -3.640 ;
        RECT 210.660 -3.980 212.960 -3.740 ;
        RECT 210.660 -4.090 211.110 -3.980 ;
        RECT 211.500 -4.420 211.910 -3.980 ;
        RECT 212.510 -4.060 212.960 -3.980 ;
        RECT 213.910 -3.740 214.360 -3.670 ;
        RECT 214.960 -3.740 215.370 -3.310 ;
        RECT 215.760 -3.740 216.210 -3.640 ;
        RECT 213.910 -3.980 216.210 -3.740 ;
        RECT 213.910 -4.090 214.360 -3.980 ;
        RECT 215.760 -4.090 216.210 -3.980 ;
        RECT 201.180 -4.640 202.710 -4.430 ;
        RECT 203.090 -4.640 203.540 -4.550 ;
        RECT 203.920 -4.640 205.450 -4.430 ;
        RECT 214.680 -4.430 215.130 -4.150 ;
        RECT 214.680 -4.640 216.210 -4.430 ;
        RECT 216.590 -4.640 217.030 -4.550 ;
        RECT 13.260 -4.900 15.370 -4.640 ;
        RECT 26.760 -4.900 28.870 -4.640 ;
        RECT 40.260 -4.900 42.370 -4.640 ;
        RECT 53.760 -4.900 55.870 -4.640 ;
        RECT 67.260 -4.900 69.370 -4.640 ;
        RECT 80.760 -4.900 82.870 -4.640 ;
        RECT 94.260 -4.900 96.370 -4.640 ;
        RECT 107.760 -4.900 109.870 -4.640 ;
        RECT 121.260 -4.900 123.370 -4.640 ;
        RECT 134.760 -4.900 136.870 -4.640 ;
        RECT 148.260 -4.900 150.370 -4.640 ;
        RECT 161.760 -4.900 163.870 -4.640 ;
        RECT 175.260 -4.900 177.370 -4.640 ;
        RECT 188.760 -4.900 190.870 -4.640 ;
        RECT 202.260 -4.900 204.370 -4.640 ;
        RECT 215.760 -4.900 217.030 -4.640 ;
        RECT 12.180 -5.110 13.710 -4.900 ;
        RECT 14.090 -4.990 14.540 -4.900 ;
        RECT 14.920 -5.110 16.450 -4.900 ;
        RECT 1.420 -5.560 1.870 -5.450 ;
        RECT 3.270 -5.560 3.720 -5.450 ;
        RECT 1.420 -5.800 3.720 -5.560 ;
        RECT 1.420 -5.900 1.870 -5.800 ;
        RECT 2.260 -6.230 2.670 -5.800 ;
        RECT 3.270 -5.870 3.720 -5.800 ;
        RECT 4.670 -5.560 5.120 -5.480 ;
        RECT 5.720 -5.560 6.130 -5.120 ;
        RECT 6.520 -5.560 6.970 -5.450 ;
        RECT 4.670 -5.800 6.970 -5.560 ;
        RECT 4.670 -5.900 5.120 -5.800 ;
        RECT 6.520 -5.900 6.970 -5.800 ;
        RECT 8.160 -5.560 8.610 -5.450 ;
        RECT 9.000 -5.560 9.410 -5.120 ;
        RECT 12.180 -5.390 12.630 -5.110 ;
        RECT 16.000 -5.390 16.450 -5.110 ;
        RECT 25.680 -5.110 27.210 -4.900 ;
        RECT 27.590 -4.990 28.040 -4.900 ;
        RECT 28.420 -5.110 29.950 -4.900 ;
        RECT 10.010 -5.560 10.460 -5.480 ;
        RECT 8.160 -5.800 10.460 -5.560 ;
        RECT 8.160 -5.900 8.610 -5.800 ;
        RECT 10.010 -5.900 10.460 -5.800 ;
        RECT 11.410 -5.560 11.860 -5.450 ;
        RECT 13.260 -5.560 13.710 -5.450 ;
        RECT 11.410 -5.800 13.710 -5.560 ;
        RECT 11.410 -5.870 11.860 -5.800 ;
        RECT 5.420 -6.380 6.970 -6.160 ;
        RECT 5.420 -6.770 5.920 -6.380 ;
        RECT 6.520 -6.430 6.970 -6.380 ;
        RECT 7.350 -6.430 7.780 -6.370 ;
        RECT 8.160 -6.380 9.710 -6.160 ;
        RECT 12.460 -6.230 12.870 -5.800 ;
        RECT 13.260 -5.900 13.710 -5.800 ;
        RECT 14.920 -5.560 15.370 -5.450 ;
        RECT 16.770 -5.560 17.220 -5.450 ;
        RECT 14.920 -5.800 17.220 -5.560 ;
        RECT 14.920 -5.900 15.370 -5.800 ;
        RECT 15.760 -6.230 16.170 -5.800 ;
        RECT 16.770 -5.870 17.220 -5.800 ;
        RECT 18.170 -5.560 18.620 -5.480 ;
        RECT 19.220 -5.560 19.630 -5.120 ;
        RECT 20.020 -5.560 20.470 -5.450 ;
        RECT 18.170 -5.800 20.470 -5.560 ;
        RECT 18.170 -5.900 18.620 -5.800 ;
        RECT 20.020 -5.900 20.470 -5.800 ;
        RECT 21.660 -5.560 22.110 -5.450 ;
        RECT 22.500 -5.560 22.910 -5.120 ;
        RECT 25.680 -5.390 26.130 -5.110 ;
        RECT 29.500 -5.390 29.950 -5.110 ;
        RECT 39.180 -5.110 40.710 -4.900 ;
        RECT 41.090 -4.990 41.540 -4.900 ;
        RECT 41.920 -5.110 43.450 -4.900 ;
        RECT 23.510 -5.560 23.960 -5.480 ;
        RECT 21.660 -5.800 23.960 -5.560 ;
        RECT 21.660 -5.900 22.110 -5.800 ;
        RECT 23.510 -5.900 23.960 -5.800 ;
        RECT 24.910 -5.560 25.360 -5.450 ;
        RECT 26.760 -5.560 27.210 -5.450 ;
        RECT 24.910 -5.800 27.210 -5.560 ;
        RECT 24.910 -5.870 25.360 -5.800 ;
        RECT 8.160 -6.430 8.610 -6.380 ;
        RECT 6.520 -6.720 8.610 -6.430 ;
        RECT 6.520 -6.770 6.970 -6.720 ;
        RECT 1.420 -7.350 1.870 -7.250 ;
        RECT 2.260 -7.350 2.670 -6.920 ;
        RECT 5.420 -6.990 6.970 -6.770 ;
        RECT 7.350 -6.780 7.780 -6.720 ;
        RECT 8.160 -6.770 8.610 -6.720 ;
        RECT 9.210 -6.770 9.710 -6.380 ;
        RECT 8.160 -6.990 9.710 -6.770 ;
        RECT 18.920 -6.380 20.470 -6.160 ;
        RECT 18.920 -6.770 19.420 -6.380 ;
        RECT 20.020 -6.430 20.470 -6.380 ;
        RECT 20.850 -6.430 21.280 -6.370 ;
        RECT 21.660 -6.380 23.210 -6.160 ;
        RECT 25.960 -6.230 26.370 -5.800 ;
        RECT 26.760 -5.900 27.210 -5.800 ;
        RECT 28.420 -5.560 28.870 -5.450 ;
        RECT 30.270 -5.560 30.720 -5.450 ;
        RECT 28.420 -5.800 30.720 -5.560 ;
        RECT 28.420 -5.900 28.870 -5.800 ;
        RECT 29.260 -6.230 29.670 -5.800 ;
        RECT 30.270 -5.870 30.720 -5.800 ;
        RECT 31.670 -5.560 32.120 -5.480 ;
        RECT 32.720 -5.560 33.130 -5.120 ;
        RECT 33.520 -5.560 33.970 -5.450 ;
        RECT 31.670 -5.800 33.970 -5.560 ;
        RECT 31.670 -5.900 32.120 -5.800 ;
        RECT 33.520 -5.900 33.970 -5.800 ;
        RECT 35.160 -5.560 35.610 -5.450 ;
        RECT 36.000 -5.560 36.410 -5.120 ;
        RECT 39.180 -5.390 39.630 -5.110 ;
        RECT 43.000 -5.390 43.450 -5.110 ;
        RECT 52.680 -5.110 54.210 -4.900 ;
        RECT 54.590 -4.990 55.040 -4.900 ;
        RECT 55.420 -5.110 56.950 -4.900 ;
        RECT 37.010 -5.560 37.460 -5.480 ;
        RECT 35.160 -5.800 37.460 -5.560 ;
        RECT 35.160 -5.900 35.610 -5.800 ;
        RECT 37.010 -5.900 37.460 -5.800 ;
        RECT 38.410 -5.560 38.860 -5.450 ;
        RECT 40.260 -5.560 40.710 -5.450 ;
        RECT 38.410 -5.800 40.710 -5.560 ;
        RECT 38.410 -5.870 38.860 -5.800 ;
        RECT 21.660 -6.430 22.110 -6.380 ;
        RECT 20.020 -6.720 22.110 -6.430 ;
        RECT 20.020 -6.770 20.470 -6.720 ;
        RECT 3.270 -7.350 3.720 -7.280 ;
        RECT 1.420 -7.590 3.720 -7.350 ;
        RECT 1.420 -7.700 1.870 -7.590 ;
        RECT 3.270 -7.700 3.720 -7.590 ;
        RECT 4.670 -7.350 5.120 -7.250 ;
        RECT 6.520 -7.350 6.970 -7.250 ;
        RECT 4.670 -7.590 6.970 -7.350 ;
        RECT 4.670 -7.670 5.120 -7.590 ;
        RECT 5.720 -8.030 6.130 -7.590 ;
        RECT 6.520 -7.700 6.970 -7.590 ;
        RECT 8.160 -7.350 8.610 -7.250 ;
        RECT 10.010 -7.350 10.460 -7.250 ;
        RECT 8.160 -7.590 10.460 -7.350 ;
        RECT 8.160 -7.700 8.610 -7.590 ;
        RECT 9.000 -8.030 9.410 -7.590 ;
        RECT 10.010 -7.670 10.460 -7.590 ;
        RECT 11.410 -7.350 11.860 -7.280 ;
        RECT 12.460 -7.350 12.870 -6.920 ;
        RECT 13.260 -7.350 13.710 -7.250 ;
        RECT 11.410 -7.590 13.710 -7.350 ;
        RECT 11.410 -7.700 11.860 -7.590 ;
        RECT 13.260 -7.700 13.710 -7.590 ;
        RECT 14.920 -7.350 15.370 -7.250 ;
        RECT 15.760 -7.350 16.170 -6.920 ;
        RECT 18.920 -6.990 20.470 -6.770 ;
        RECT 20.850 -6.780 21.280 -6.720 ;
        RECT 21.660 -6.770 22.110 -6.720 ;
        RECT 22.710 -6.770 23.210 -6.380 ;
        RECT 21.660 -6.990 23.210 -6.770 ;
        RECT 32.420 -6.380 33.970 -6.160 ;
        RECT 32.420 -6.770 32.920 -6.380 ;
        RECT 33.520 -6.430 33.970 -6.380 ;
        RECT 34.350 -6.430 34.780 -6.370 ;
        RECT 35.160 -6.380 36.710 -6.160 ;
        RECT 39.460 -6.230 39.870 -5.800 ;
        RECT 40.260 -5.900 40.710 -5.800 ;
        RECT 41.920 -5.560 42.370 -5.450 ;
        RECT 43.770 -5.560 44.220 -5.450 ;
        RECT 41.920 -5.800 44.220 -5.560 ;
        RECT 41.920 -5.900 42.370 -5.800 ;
        RECT 42.760 -6.230 43.170 -5.800 ;
        RECT 43.770 -5.870 44.220 -5.800 ;
        RECT 45.170 -5.560 45.620 -5.480 ;
        RECT 46.220 -5.560 46.630 -5.120 ;
        RECT 47.020 -5.560 47.470 -5.450 ;
        RECT 45.170 -5.800 47.470 -5.560 ;
        RECT 45.170 -5.900 45.620 -5.800 ;
        RECT 47.020 -5.900 47.470 -5.800 ;
        RECT 48.660 -5.560 49.110 -5.450 ;
        RECT 49.500 -5.560 49.910 -5.120 ;
        RECT 52.680 -5.390 53.130 -5.110 ;
        RECT 56.500 -5.390 56.950 -5.110 ;
        RECT 66.180 -5.110 67.710 -4.900 ;
        RECT 68.090 -4.990 68.540 -4.900 ;
        RECT 68.920 -5.110 70.450 -4.900 ;
        RECT 50.510 -5.560 50.960 -5.480 ;
        RECT 48.660 -5.800 50.960 -5.560 ;
        RECT 48.660 -5.900 49.110 -5.800 ;
        RECT 50.510 -5.900 50.960 -5.800 ;
        RECT 51.910 -5.560 52.360 -5.450 ;
        RECT 53.760 -5.560 54.210 -5.450 ;
        RECT 51.910 -5.800 54.210 -5.560 ;
        RECT 51.910 -5.870 52.360 -5.800 ;
        RECT 35.160 -6.430 35.610 -6.380 ;
        RECT 33.520 -6.720 35.610 -6.430 ;
        RECT 33.520 -6.770 33.970 -6.720 ;
        RECT 16.770 -7.350 17.220 -7.280 ;
        RECT 14.920 -7.590 17.220 -7.350 ;
        RECT 14.920 -7.700 15.370 -7.590 ;
        RECT 16.770 -7.700 17.220 -7.590 ;
        RECT 18.170 -7.350 18.620 -7.250 ;
        RECT 20.020 -7.350 20.470 -7.250 ;
        RECT 18.170 -7.590 20.470 -7.350 ;
        RECT 18.170 -7.670 18.620 -7.590 ;
        RECT 12.180 -8.040 12.630 -7.760 ;
        RECT 16.000 -8.040 16.450 -7.760 ;
        RECT 19.220 -8.030 19.630 -7.590 ;
        RECT 20.020 -7.700 20.470 -7.590 ;
        RECT 21.660 -7.350 22.110 -7.250 ;
        RECT 23.510 -7.350 23.960 -7.250 ;
        RECT 21.660 -7.590 23.960 -7.350 ;
        RECT 21.660 -7.700 22.110 -7.590 ;
        RECT 22.500 -8.030 22.910 -7.590 ;
        RECT 23.510 -7.670 23.960 -7.590 ;
        RECT 24.910 -7.350 25.360 -7.280 ;
        RECT 25.960 -7.350 26.370 -6.920 ;
        RECT 26.760 -7.350 27.210 -7.250 ;
        RECT 24.910 -7.590 27.210 -7.350 ;
        RECT 24.910 -7.700 25.360 -7.590 ;
        RECT 26.760 -7.700 27.210 -7.590 ;
        RECT 28.420 -7.350 28.870 -7.250 ;
        RECT 29.260 -7.350 29.670 -6.920 ;
        RECT 32.420 -6.990 33.970 -6.770 ;
        RECT 34.350 -6.780 34.780 -6.720 ;
        RECT 35.160 -6.770 35.610 -6.720 ;
        RECT 36.210 -6.770 36.710 -6.380 ;
        RECT 35.160 -6.990 36.710 -6.770 ;
        RECT 45.920 -6.380 47.470 -6.160 ;
        RECT 45.920 -6.770 46.420 -6.380 ;
        RECT 47.020 -6.430 47.470 -6.380 ;
        RECT 47.850 -6.430 48.280 -6.370 ;
        RECT 48.660 -6.380 50.210 -6.160 ;
        RECT 52.960 -6.230 53.370 -5.800 ;
        RECT 53.760 -5.900 54.210 -5.800 ;
        RECT 55.420 -5.560 55.870 -5.450 ;
        RECT 57.270 -5.560 57.720 -5.450 ;
        RECT 55.420 -5.800 57.720 -5.560 ;
        RECT 55.420 -5.900 55.870 -5.800 ;
        RECT 56.260 -6.230 56.670 -5.800 ;
        RECT 57.270 -5.870 57.720 -5.800 ;
        RECT 58.670 -5.560 59.120 -5.480 ;
        RECT 59.720 -5.560 60.130 -5.120 ;
        RECT 60.520 -5.560 60.970 -5.450 ;
        RECT 58.670 -5.800 60.970 -5.560 ;
        RECT 58.670 -5.900 59.120 -5.800 ;
        RECT 60.520 -5.900 60.970 -5.800 ;
        RECT 62.160 -5.560 62.610 -5.450 ;
        RECT 63.000 -5.560 63.410 -5.120 ;
        RECT 66.180 -5.390 66.630 -5.110 ;
        RECT 70.000 -5.390 70.450 -5.110 ;
        RECT 79.680 -5.110 81.210 -4.900 ;
        RECT 81.590 -4.990 82.040 -4.900 ;
        RECT 82.420 -5.110 83.950 -4.900 ;
        RECT 64.010 -5.560 64.460 -5.480 ;
        RECT 62.160 -5.800 64.460 -5.560 ;
        RECT 62.160 -5.900 62.610 -5.800 ;
        RECT 64.010 -5.900 64.460 -5.800 ;
        RECT 65.410 -5.560 65.860 -5.450 ;
        RECT 67.260 -5.560 67.710 -5.450 ;
        RECT 65.410 -5.800 67.710 -5.560 ;
        RECT 65.410 -5.870 65.860 -5.800 ;
        RECT 48.660 -6.430 49.110 -6.380 ;
        RECT 47.020 -6.720 49.110 -6.430 ;
        RECT 47.020 -6.770 47.470 -6.720 ;
        RECT 30.270 -7.350 30.720 -7.280 ;
        RECT 28.420 -7.590 30.720 -7.350 ;
        RECT 28.420 -7.700 28.870 -7.590 ;
        RECT 30.270 -7.700 30.720 -7.590 ;
        RECT 31.670 -7.350 32.120 -7.250 ;
        RECT 33.520 -7.350 33.970 -7.250 ;
        RECT 31.670 -7.590 33.970 -7.350 ;
        RECT 31.670 -7.670 32.120 -7.590 ;
        RECT 12.180 -8.250 13.710 -8.040 ;
        RECT 14.090 -8.250 14.540 -8.160 ;
        RECT 14.920 -8.250 16.450 -8.040 ;
        RECT 25.680 -8.040 26.130 -7.760 ;
        RECT 29.500 -8.040 29.950 -7.760 ;
        RECT 32.720 -8.030 33.130 -7.590 ;
        RECT 33.520 -7.700 33.970 -7.590 ;
        RECT 35.160 -7.350 35.610 -7.250 ;
        RECT 37.010 -7.350 37.460 -7.250 ;
        RECT 35.160 -7.590 37.460 -7.350 ;
        RECT 35.160 -7.700 35.610 -7.590 ;
        RECT 36.000 -8.030 36.410 -7.590 ;
        RECT 37.010 -7.670 37.460 -7.590 ;
        RECT 38.410 -7.350 38.860 -7.280 ;
        RECT 39.460 -7.350 39.870 -6.920 ;
        RECT 40.260 -7.350 40.710 -7.250 ;
        RECT 38.410 -7.590 40.710 -7.350 ;
        RECT 38.410 -7.700 38.860 -7.590 ;
        RECT 40.260 -7.700 40.710 -7.590 ;
        RECT 41.920 -7.350 42.370 -7.250 ;
        RECT 42.760 -7.350 43.170 -6.920 ;
        RECT 45.920 -6.990 47.470 -6.770 ;
        RECT 47.850 -6.780 48.280 -6.720 ;
        RECT 48.660 -6.770 49.110 -6.720 ;
        RECT 49.710 -6.770 50.210 -6.380 ;
        RECT 48.660 -6.990 50.210 -6.770 ;
        RECT 59.420 -6.380 60.970 -6.160 ;
        RECT 59.420 -6.770 59.920 -6.380 ;
        RECT 60.520 -6.430 60.970 -6.380 ;
        RECT 61.350 -6.430 61.780 -6.370 ;
        RECT 62.160 -6.380 63.710 -6.160 ;
        RECT 66.460 -6.230 66.870 -5.800 ;
        RECT 67.260 -5.900 67.710 -5.800 ;
        RECT 68.920 -5.560 69.370 -5.450 ;
        RECT 70.770 -5.560 71.220 -5.450 ;
        RECT 68.920 -5.800 71.220 -5.560 ;
        RECT 68.920 -5.900 69.370 -5.800 ;
        RECT 69.760 -6.230 70.170 -5.800 ;
        RECT 70.770 -5.870 71.220 -5.800 ;
        RECT 72.170 -5.560 72.620 -5.480 ;
        RECT 73.220 -5.560 73.630 -5.120 ;
        RECT 74.020 -5.560 74.470 -5.450 ;
        RECT 72.170 -5.800 74.470 -5.560 ;
        RECT 72.170 -5.900 72.620 -5.800 ;
        RECT 74.020 -5.900 74.470 -5.800 ;
        RECT 75.660 -5.560 76.110 -5.450 ;
        RECT 76.500 -5.560 76.910 -5.120 ;
        RECT 79.680 -5.390 80.130 -5.110 ;
        RECT 83.500 -5.390 83.950 -5.110 ;
        RECT 93.180 -5.110 94.710 -4.900 ;
        RECT 95.090 -4.990 95.540 -4.900 ;
        RECT 95.920 -5.110 97.450 -4.900 ;
        RECT 77.510 -5.560 77.960 -5.480 ;
        RECT 75.660 -5.800 77.960 -5.560 ;
        RECT 75.660 -5.900 76.110 -5.800 ;
        RECT 77.510 -5.900 77.960 -5.800 ;
        RECT 78.910 -5.560 79.360 -5.450 ;
        RECT 80.760 -5.560 81.210 -5.450 ;
        RECT 78.910 -5.800 81.210 -5.560 ;
        RECT 78.910 -5.870 79.360 -5.800 ;
        RECT 62.160 -6.430 62.610 -6.380 ;
        RECT 60.520 -6.720 62.610 -6.430 ;
        RECT 60.520 -6.770 60.970 -6.720 ;
        RECT 43.770 -7.350 44.220 -7.280 ;
        RECT 41.920 -7.590 44.220 -7.350 ;
        RECT 41.920 -7.700 42.370 -7.590 ;
        RECT 43.770 -7.700 44.220 -7.590 ;
        RECT 45.170 -7.350 45.620 -7.250 ;
        RECT 47.020 -7.350 47.470 -7.250 ;
        RECT 45.170 -7.590 47.470 -7.350 ;
        RECT 45.170 -7.670 45.620 -7.590 ;
        RECT 25.680 -8.250 27.210 -8.040 ;
        RECT 27.590 -8.250 28.040 -8.160 ;
        RECT 28.420 -8.250 29.950 -8.040 ;
        RECT 39.180 -8.040 39.630 -7.760 ;
        RECT 43.000 -8.040 43.450 -7.760 ;
        RECT 46.220 -8.030 46.630 -7.590 ;
        RECT 47.020 -7.700 47.470 -7.590 ;
        RECT 48.660 -7.350 49.110 -7.250 ;
        RECT 50.510 -7.350 50.960 -7.250 ;
        RECT 48.660 -7.590 50.960 -7.350 ;
        RECT 48.660 -7.700 49.110 -7.590 ;
        RECT 49.500 -8.030 49.910 -7.590 ;
        RECT 50.510 -7.670 50.960 -7.590 ;
        RECT 51.910 -7.350 52.360 -7.280 ;
        RECT 52.960 -7.350 53.370 -6.920 ;
        RECT 53.760 -7.350 54.210 -7.250 ;
        RECT 51.910 -7.590 54.210 -7.350 ;
        RECT 51.910 -7.700 52.360 -7.590 ;
        RECT 53.760 -7.700 54.210 -7.590 ;
        RECT 55.420 -7.350 55.870 -7.250 ;
        RECT 56.260 -7.350 56.670 -6.920 ;
        RECT 59.420 -6.990 60.970 -6.770 ;
        RECT 61.350 -6.780 61.780 -6.720 ;
        RECT 62.160 -6.770 62.610 -6.720 ;
        RECT 63.210 -6.770 63.710 -6.380 ;
        RECT 62.160 -6.990 63.710 -6.770 ;
        RECT 72.920 -6.380 74.470 -6.160 ;
        RECT 72.920 -6.770 73.420 -6.380 ;
        RECT 74.020 -6.430 74.470 -6.380 ;
        RECT 74.850 -6.430 75.280 -6.370 ;
        RECT 75.660 -6.380 77.210 -6.160 ;
        RECT 79.960 -6.230 80.370 -5.800 ;
        RECT 80.760 -5.900 81.210 -5.800 ;
        RECT 82.420 -5.560 82.870 -5.450 ;
        RECT 84.270 -5.560 84.720 -5.450 ;
        RECT 82.420 -5.800 84.720 -5.560 ;
        RECT 82.420 -5.900 82.870 -5.800 ;
        RECT 83.260 -6.230 83.670 -5.800 ;
        RECT 84.270 -5.870 84.720 -5.800 ;
        RECT 85.670 -5.560 86.120 -5.480 ;
        RECT 86.720 -5.560 87.130 -5.120 ;
        RECT 87.520 -5.560 87.970 -5.450 ;
        RECT 85.670 -5.800 87.970 -5.560 ;
        RECT 85.670 -5.900 86.120 -5.800 ;
        RECT 87.520 -5.900 87.970 -5.800 ;
        RECT 89.160 -5.560 89.610 -5.450 ;
        RECT 90.000 -5.560 90.410 -5.120 ;
        RECT 93.180 -5.390 93.630 -5.110 ;
        RECT 97.000 -5.390 97.450 -5.110 ;
        RECT 106.680 -5.110 108.210 -4.900 ;
        RECT 108.590 -4.990 109.040 -4.900 ;
        RECT 109.420 -5.110 110.950 -4.900 ;
        RECT 91.010 -5.560 91.460 -5.480 ;
        RECT 89.160 -5.800 91.460 -5.560 ;
        RECT 89.160 -5.900 89.610 -5.800 ;
        RECT 91.010 -5.900 91.460 -5.800 ;
        RECT 92.410 -5.560 92.860 -5.450 ;
        RECT 94.260 -5.560 94.710 -5.450 ;
        RECT 92.410 -5.800 94.710 -5.560 ;
        RECT 92.410 -5.870 92.860 -5.800 ;
        RECT 75.660 -6.430 76.110 -6.380 ;
        RECT 74.020 -6.720 76.110 -6.430 ;
        RECT 74.020 -6.770 74.470 -6.720 ;
        RECT 57.270 -7.350 57.720 -7.280 ;
        RECT 55.420 -7.590 57.720 -7.350 ;
        RECT 55.420 -7.700 55.870 -7.590 ;
        RECT 57.270 -7.700 57.720 -7.590 ;
        RECT 58.670 -7.350 59.120 -7.250 ;
        RECT 60.520 -7.350 60.970 -7.250 ;
        RECT 58.670 -7.590 60.970 -7.350 ;
        RECT 58.670 -7.670 59.120 -7.590 ;
        RECT 39.180 -8.250 40.710 -8.040 ;
        RECT 41.090 -8.250 41.540 -8.160 ;
        RECT 41.920 -8.250 43.450 -8.040 ;
        RECT 52.680 -8.040 53.130 -7.760 ;
        RECT 56.500 -8.040 56.950 -7.760 ;
        RECT 59.720 -8.030 60.130 -7.590 ;
        RECT 60.520 -7.700 60.970 -7.590 ;
        RECT 62.160 -7.350 62.610 -7.250 ;
        RECT 64.010 -7.350 64.460 -7.250 ;
        RECT 62.160 -7.590 64.460 -7.350 ;
        RECT 62.160 -7.700 62.610 -7.590 ;
        RECT 63.000 -8.030 63.410 -7.590 ;
        RECT 64.010 -7.670 64.460 -7.590 ;
        RECT 65.410 -7.350 65.860 -7.280 ;
        RECT 66.460 -7.350 66.870 -6.920 ;
        RECT 67.260 -7.350 67.710 -7.250 ;
        RECT 65.410 -7.590 67.710 -7.350 ;
        RECT 65.410 -7.700 65.860 -7.590 ;
        RECT 67.260 -7.700 67.710 -7.590 ;
        RECT 68.920 -7.350 69.370 -7.250 ;
        RECT 69.760 -7.350 70.170 -6.920 ;
        RECT 72.920 -6.990 74.470 -6.770 ;
        RECT 74.850 -6.780 75.280 -6.720 ;
        RECT 75.660 -6.770 76.110 -6.720 ;
        RECT 76.710 -6.770 77.210 -6.380 ;
        RECT 75.660 -6.990 77.210 -6.770 ;
        RECT 86.420 -6.380 87.970 -6.160 ;
        RECT 86.420 -6.770 86.920 -6.380 ;
        RECT 87.520 -6.430 87.970 -6.380 ;
        RECT 88.350 -6.430 88.780 -6.370 ;
        RECT 89.160 -6.380 90.710 -6.160 ;
        RECT 93.460 -6.230 93.870 -5.800 ;
        RECT 94.260 -5.900 94.710 -5.800 ;
        RECT 95.920 -5.560 96.370 -5.450 ;
        RECT 97.770 -5.560 98.220 -5.450 ;
        RECT 95.920 -5.800 98.220 -5.560 ;
        RECT 95.920 -5.900 96.370 -5.800 ;
        RECT 96.760 -6.230 97.170 -5.800 ;
        RECT 97.770 -5.870 98.220 -5.800 ;
        RECT 99.170 -5.560 99.620 -5.480 ;
        RECT 100.220 -5.560 100.630 -5.120 ;
        RECT 101.020 -5.560 101.470 -5.450 ;
        RECT 99.170 -5.800 101.470 -5.560 ;
        RECT 99.170 -5.900 99.620 -5.800 ;
        RECT 101.020 -5.900 101.470 -5.800 ;
        RECT 102.660 -5.560 103.110 -5.450 ;
        RECT 103.500 -5.560 103.910 -5.120 ;
        RECT 106.680 -5.390 107.130 -5.110 ;
        RECT 110.500 -5.390 110.950 -5.110 ;
        RECT 120.180 -5.110 121.710 -4.900 ;
        RECT 122.090 -4.990 122.540 -4.900 ;
        RECT 122.920 -5.110 124.450 -4.900 ;
        RECT 104.510 -5.560 104.960 -5.480 ;
        RECT 102.660 -5.800 104.960 -5.560 ;
        RECT 102.660 -5.900 103.110 -5.800 ;
        RECT 104.510 -5.900 104.960 -5.800 ;
        RECT 105.910 -5.560 106.360 -5.450 ;
        RECT 107.760 -5.560 108.210 -5.450 ;
        RECT 105.910 -5.800 108.210 -5.560 ;
        RECT 105.910 -5.870 106.360 -5.800 ;
        RECT 89.160 -6.430 89.610 -6.380 ;
        RECT 87.520 -6.720 89.610 -6.430 ;
        RECT 87.520 -6.770 87.970 -6.720 ;
        RECT 70.770 -7.350 71.220 -7.280 ;
        RECT 68.920 -7.590 71.220 -7.350 ;
        RECT 68.920 -7.700 69.370 -7.590 ;
        RECT 70.770 -7.700 71.220 -7.590 ;
        RECT 72.170 -7.350 72.620 -7.250 ;
        RECT 74.020 -7.350 74.470 -7.250 ;
        RECT 72.170 -7.590 74.470 -7.350 ;
        RECT 72.170 -7.670 72.620 -7.590 ;
        RECT 52.680 -8.250 54.210 -8.040 ;
        RECT 54.590 -8.250 55.040 -8.160 ;
        RECT 55.420 -8.250 56.950 -8.040 ;
        RECT 66.180 -8.040 66.630 -7.760 ;
        RECT 70.000 -8.040 70.450 -7.760 ;
        RECT 73.220 -8.030 73.630 -7.590 ;
        RECT 74.020 -7.700 74.470 -7.590 ;
        RECT 75.660 -7.350 76.110 -7.250 ;
        RECT 77.510 -7.350 77.960 -7.250 ;
        RECT 75.660 -7.590 77.960 -7.350 ;
        RECT 75.660 -7.700 76.110 -7.590 ;
        RECT 76.500 -8.030 76.910 -7.590 ;
        RECT 77.510 -7.670 77.960 -7.590 ;
        RECT 78.910 -7.350 79.360 -7.280 ;
        RECT 79.960 -7.350 80.370 -6.920 ;
        RECT 80.760 -7.350 81.210 -7.250 ;
        RECT 78.910 -7.590 81.210 -7.350 ;
        RECT 78.910 -7.700 79.360 -7.590 ;
        RECT 80.760 -7.700 81.210 -7.590 ;
        RECT 82.420 -7.350 82.870 -7.250 ;
        RECT 83.260 -7.350 83.670 -6.920 ;
        RECT 86.420 -6.990 87.970 -6.770 ;
        RECT 88.350 -6.780 88.780 -6.720 ;
        RECT 89.160 -6.770 89.610 -6.720 ;
        RECT 90.210 -6.770 90.710 -6.380 ;
        RECT 89.160 -6.990 90.710 -6.770 ;
        RECT 99.920 -6.380 101.470 -6.160 ;
        RECT 99.920 -6.770 100.420 -6.380 ;
        RECT 101.020 -6.430 101.470 -6.380 ;
        RECT 101.850 -6.430 102.280 -6.370 ;
        RECT 102.660 -6.380 104.210 -6.160 ;
        RECT 106.960 -6.230 107.370 -5.800 ;
        RECT 107.760 -5.900 108.210 -5.800 ;
        RECT 109.420 -5.560 109.870 -5.450 ;
        RECT 111.270 -5.560 111.720 -5.450 ;
        RECT 109.420 -5.800 111.720 -5.560 ;
        RECT 109.420 -5.900 109.870 -5.800 ;
        RECT 110.260 -6.230 110.670 -5.800 ;
        RECT 111.270 -5.870 111.720 -5.800 ;
        RECT 112.670 -5.560 113.120 -5.480 ;
        RECT 113.720 -5.560 114.130 -5.120 ;
        RECT 114.520 -5.560 114.970 -5.450 ;
        RECT 112.670 -5.800 114.970 -5.560 ;
        RECT 112.670 -5.900 113.120 -5.800 ;
        RECT 114.520 -5.900 114.970 -5.800 ;
        RECT 116.160 -5.560 116.610 -5.450 ;
        RECT 117.000 -5.560 117.410 -5.120 ;
        RECT 120.180 -5.390 120.630 -5.110 ;
        RECT 124.000 -5.390 124.450 -5.110 ;
        RECT 133.680 -5.110 135.210 -4.900 ;
        RECT 135.590 -4.990 136.040 -4.900 ;
        RECT 136.420 -5.110 137.950 -4.900 ;
        RECT 118.010 -5.560 118.460 -5.480 ;
        RECT 116.160 -5.800 118.460 -5.560 ;
        RECT 116.160 -5.900 116.610 -5.800 ;
        RECT 118.010 -5.900 118.460 -5.800 ;
        RECT 119.410 -5.560 119.860 -5.450 ;
        RECT 121.260 -5.560 121.710 -5.450 ;
        RECT 119.410 -5.800 121.710 -5.560 ;
        RECT 119.410 -5.870 119.860 -5.800 ;
        RECT 102.660 -6.430 103.110 -6.380 ;
        RECT 101.020 -6.720 103.110 -6.430 ;
        RECT 101.020 -6.770 101.470 -6.720 ;
        RECT 84.270 -7.350 84.720 -7.280 ;
        RECT 82.420 -7.590 84.720 -7.350 ;
        RECT 82.420 -7.700 82.870 -7.590 ;
        RECT 84.270 -7.700 84.720 -7.590 ;
        RECT 85.670 -7.350 86.120 -7.250 ;
        RECT 87.520 -7.350 87.970 -7.250 ;
        RECT 85.670 -7.590 87.970 -7.350 ;
        RECT 85.670 -7.670 86.120 -7.590 ;
        RECT 66.180 -8.250 67.710 -8.040 ;
        RECT 68.090 -8.250 68.540 -8.160 ;
        RECT 68.920 -8.250 70.450 -8.040 ;
        RECT 79.680 -8.040 80.130 -7.760 ;
        RECT 83.500 -8.040 83.950 -7.760 ;
        RECT 86.720 -8.030 87.130 -7.590 ;
        RECT 87.520 -7.700 87.970 -7.590 ;
        RECT 89.160 -7.350 89.610 -7.250 ;
        RECT 91.010 -7.350 91.460 -7.250 ;
        RECT 89.160 -7.590 91.460 -7.350 ;
        RECT 89.160 -7.700 89.610 -7.590 ;
        RECT 90.000 -8.030 90.410 -7.590 ;
        RECT 91.010 -7.670 91.460 -7.590 ;
        RECT 92.410 -7.350 92.860 -7.280 ;
        RECT 93.460 -7.350 93.870 -6.920 ;
        RECT 94.260 -7.350 94.710 -7.250 ;
        RECT 92.410 -7.590 94.710 -7.350 ;
        RECT 92.410 -7.700 92.860 -7.590 ;
        RECT 94.260 -7.700 94.710 -7.590 ;
        RECT 95.920 -7.350 96.370 -7.250 ;
        RECT 96.760 -7.350 97.170 -6.920 ;
        RECT 99.920 -6.990 101.470 -6.770 ;
        RECT 101.850 -6.780 102.280 -6.720 ;
        RECT 102.660 -6.770 103.110 -6.720 ;
        RECT 103.710 -6.770 104.210 -6.380 ;
        RECT 102.660 -6.990 104.210 -6.770 ;
        RECT 113.420 -6.380 114.970 -6.160 ;
        RECT 113.420 -6.770 113.920 -6.380 ;
        RECT 114.520 -6.430 114.970 -6.380 ;
        RECT 115.350 -6.430 115.780 -6.370 ;
        RECT 116.160 -6.380 117.710 -6.160 ;
        RECT 120.460 -6.230 120.870 -5.800 ;
        RECT 121.260 -5.900 121.710 -5.800 ;
        RECT 122.920 -5.560 123.370 -5.450 ;
        RECT 124.770 -5.560 125.220 -5.450 ;
        RECT 122.920 -5.800 125.220 -5.560 ;
        RECT 122.920 -5.900 123.370 -5.800 ;
        RECT 123.760 -6.230 124.170 -5.800 ;
        RECT 124.770 -5.870 125.220 -5.800 ;
        RECT 126.170 -5.560 126.620 -5.480 ;
        RECT 127.220 -5.560 127.630 -5.120 ;
        RECT 128.020 -5.560 128.470 -5.450 ;
        RECT 126.170 -5.800 128.470 -5.560 ;
        RECT 126.170 -5.900 126.620 -5.800 ;
        RECT 128.020 -5.900 128.470 -5.800 ;
        RECT 129.660 -5.560 130.110 -5.450 ;
        RECT 130.500 -5.560 130.910 -5.120 ;
        RECT 133.680 -5.390 134.130 -5.110 ;
        RECT 137.500 -5.390 137.950 -5.110 ;
        RECT 147.180 -5.110 148.710 -4.900 ;
        RECT 149.090 -4.990 149.540 -4.900 ;
        RECT 149.920 -5.110 151.450 -4.900 ;
        RECT 131.510 -5.560 131.960 -5.480 ;
        RECT 129.660 -5.800 131.960 -5.560 ;
        RECT 129.660 -5.900 130.110 -5.800 ;
        RECT 131.510 -5.900 131.960 -5.800 ;
        RECT 132.910 -5.560 133.360 -5.450 ;
        RECT 134.760 -5.560 135.210 -5.450 ;
        RECT 132.910 -5.800 135.210 -5.560 ;
        RECT 132.910 -5.870 133.360 -5.800 ;
        RECT 116.160 -6.430 116.610 -6.380 ;
        RECT 114.520 -6.720 116.610 -6.430 ;
        RECT 114.520 -6.770 114.970 -6.720 ;
        RECT 97.770 -7.350 98.220 -7.280 ;
        RECT 95.920 -7.590 98.220 -7.350 ;
        RECT 95.920 -7.700 96.370 -7.590 ;
        RECT 97.770 -7.700 98.220 -7.590 ;
        RECT 99.170 -7.350 99.620 -7.250 ;
        RECT 101.020 -7.350 101.470 -7.250 ;
        RECT 99.170 -7.590 101.470 -7.350 ;
        RECT 99.170 -7.670 99.620 -7.590 ;
        RECT 79.680 -8.250 81.210 -8.040 ;
        RECT 81.590 -8.250 82.040 -8.160 ;
        RECT 82.420 -8.250 83.950 -8.040 ;
        RECT 93.180 -8.040 93.630 -7.760 ;
        RECT 97.000 -8.040 97.450 -7.760 ;
        RECT 100.220 -8.030 100.630 -7.590 ;
        RECT 101.020 -7.700 101.470 -7.590 ;
        RECT 102.660 -7.350 103.110 -7.250 ;
        RECT 104.510 -7.350 104.960 -7.250 ;
        RECT 102.660 -7.590 104.960 -7.350 ;
        RECT 102.660 -7.700 103.110 -7.590 ;
        RECT 103.500 -8.030 103.910 -7.590 ;
        RECT 104.510 -7.670 104.960 -7.590 ;
        RECT 105.910 -7.350 106.360 -7.280 ;
        RECT 106.960 -7.350 107.370 -6.920 ;
        RECT 107.760 -7.350 108.210 -7.250 ;
        RECT 105.910 -7.590 108.210 -7.350 ;
        RECT 105.910 -7.700 106.360 -7.590 ;
        RECT 107.760 -7.700 108.210 -7.590 ;
        RECT 109.420 -7.350 109.870 -7.250 ;
        RECT 110.260 -7.350 110.670 -6.920 ;
        RECT 113.420 -6.990 114.970 -6.770 ;
        RECT 115.350 -6.780 115.780 -6.720 ;
        RECT 116.160 -6.770 116.610 -6.720 ;
        RECT 117.210 -6.770 117.710 -6.380 ;
        RECT 116.160 -6.990 117.710 -6.770 ;
        RECT 126.920 -6.380 128.470 -6.160 ;
        RECT 126.920 -6.770 127.420 -6.380 ;
        RECT 128.020 -6.430 128.470 -6.380 ;
        RECT 128.850 -6.430 129.280 -6.370 ;
        RECT 129.660 -6.380 131.210 -6.160 ;
        RECT 133.960 -6.230 134.370 -5.800 ;
        RECT 134.760 -5.900 135.210 -5.800 ;
        RECT 136.420 -5.560 136.870 -5.450 ;
        RECT 138.270 -5.560 138.720 -5.450 ;
        RECT 136.420 -5.800 138.720 -5.560 ;
        RECT 136.420 -5.900 136.870 -5.800 ;
        RECT 137.260 -6.230 137.670 -5.800 ;
        RECT 138.270 -5.870 138.720 -5.800 ;
        RECT 139.670 -5.560 140.120 -5.480 ;
        RECT 140.720 -5.560 141.130 -5.120 ;
        RECT 141.520 -5.560 141.970 -5.450 ;
        RECT 139.670 -5.800 141.970 -5.560 ;
        RECT 139.670 -5.900 140.120 -5.800 ;
        RECT 141.520 -5.900 141.970 -5.800 ;
        RECT 143.160 -5.560 143.610 -5.450 ;
        RECT 144.000 -5.560 144.410 -5.120 ;
        RECT 147.180 -5.390 147.630 -5.110 ;
        RECT 151.000 -5.390 151.450 -5.110 ;
        RECT 160.680 -5.110 162.210 -4.900 ;
        RECT 162.590 -4.990 163.040 -4.900 ;
        RECT 163.420 -5.110 164.950 -4.900 ;
        RECT 145.010 -5.560 145.460 -5.480 ;
        RECT 143.160 -5.800 145.460 -5.560 ;
        RECT 143.160 -5.900 143.610 -5.800 ;
        RECT 145.010 -5.900 145.460 -5.800 ;
        RECT 146.410 -5.560 146.860 -5.450 ;
        RECT 148.260 -5.560 148.710 -5.450 ;
        RECT 146.410 -5.800 148.710 -5.560 ;
        RECT 146.410 -5.870 146.860 -5.800 ;
        RECT 129.660 -6.430 130.110 -6.380 ;
        RECT 128.020 -6.720 130.110 -6.430 ;
        RECT 128.020 -6.770 128.470 -6.720 ;
        RECT 111.270 -7.350 111.720 -7.280 ;
        RECT 109.420 -7.590 111.720 -7.350 ;
        RECT 109.420 -7.700 109.870 -7.590 ;
        RECT 111.270 -7.700 111.720 -7.590 ;
        RECT 112.670 -7.350 113.120 -7.250 ;
        RECT 114.520 -7.350 114.970 -7.250 ;
        RECT 112.670 -7.590 114.970 -7.350 ;
        RECT 112.670 -7.670 113.120 -7.590 ;
        RECT 93.180 -8.250 94.710 -8.040 ;
        RECT 95.090 -8.250 95.540 -8.160 ;
        RECT 95.920 -8.250 97.450 -8.040 ;
        RECT 106.680 -8.040 107.130 -7.760 ;
        RECT 110.500 -8.040 110.950 -7.760 ;
        RECT 113.720 -8.030 114.130 -7.590 ;
        RECT 114.520 -7.700 114.970 -7.590 ;
        RECT 116.160 -7.350 116.610 -7.250 ;
        RECT 118.010 -7.350 118.460 -7.250 ;
        RECT 116.160 -7.590 118.460 -7.350 ;
        RECT 116.160 -7.700 116.610 -7.590 ;
        RECT 117.000 -8.030 117.410 -7.590 ;
        RECT 118.010 -7.670 118.460 -7.590 ;
        RECT 119.410 -7.350 119.860 -7.280 ;
        RECT 120.460 -7.350 120.870 -6.920 ;
        RECT 121.260 -7.350 121.710 -7.250 ;
        RECT 119.410 -7.590 121.710 -7.350 ;
        RECT 119.410 -7.700 119.860 -7.590 ;
        RECT 121.260 -7.700 121.710 -7.590 ;
        RECT 122.920 -7.350 123.370 -7.250 ;
        RECT 123.760 -7.350 124.170 -6.920 ;
        RECT 126.920 -6.990 128.470 -6.770 ;
        RECT 128.850 -6.780 129.280 -6.720 ;
        RECT 129.660 -6.770 130.110 -6.720 ;
        RECT 130.710 -6.770 131.210 -6.380 ;
        RECT 129.660 -6.990 131.210 -6.770 ;
        RECT 140.420 -6.380 141.970 -6.160 ;
        RECT 140.420 -6.770 140.920 -6.380 ;
        RECT 141.520 -6.430 141.970 -6.380 ;
        RECT 142.350 -6.430 142.780 -6.370 ;
        RECT 143.160 -6.380 144.710 -6.160 ;
        RECT 147.460 -6.230 147.870 -5.800 ;
        RECT 148.260 -5.900 148.710 -5.800 ;
        RECT 149.920 -5.560 150.370 -5.450 ;
        RECT 151.770 -5.560 152.220 -5.450 ;
        RECT 149.920 -5.800 152.220 -5.560 ;
        RECT 149.920 -5.900 150.370 -5.800 ;
        RECT 150.760 -6.230 151.170 -5.800 ;
        RECT 151.770 -5.870 152.220 -5.800 ;
        RECT 153.170 -5.560 153.620 -5.480 ;
        RECT 154.220 -5.560 154.630 -5.120 ;
        RECT 155.020 -5.560 155.470 -5.450 ;
        RECT 153.170 -5.800 155.470 -5.560 ;
        RECT 153.170 -5.900 153.620 -5.800 ;
        RECT 155.020 -5.900 155.470 -5.800 ;
        RECT 156.660 -5.560 157.110 -5.450 ;
        RECT 157.500 -5.560 157.910 -5.120 ;
        RECT 160.680 -5.390 161.130 -5.110 ;
        RECT 164.500 -5.390 164.950 -5.110 ;
        RECT 174.180 -5.110 175.710 -4.900 ;
        RECT 176.090 -4.990 176.540 -4.900 ;
        RECT 176.920 -5.110 178.450 -4.900 ;
        RECT 158.510 -5.560 158.960 -5.480 ;
        RECT 156.660 -5.800 158.960 -5.560 ;
        RECT 156.660 -5.900 157.110 -5.800 ;
        RECT 158.510 -5.900 158.960 -5.800 ;
        RECT 159.910 -5.560 160.360 -5.450 ;
        RECT 161.760 -5.560 162.210 -5.450 ;
        RECT 159.910 -5.800 162.210 -5.560 ;
        RECT 159.910 -5.870 160.360 -5.800 ;
        RECT 143.160 -6.430 143.610 -6.380 ;
        RECT 141.520 -6.720 143.610 -6.430 ;
        RECT 141.520 -6.770 141.970 -6.720 ;
        RECT 124.770 -7.350 125.220 -7.280 ;
        RECT 122.920 -7.590 125.220 -7.350 ;
        RECT 122.920 -7.700 123.370 -7.590 ;
        RECT 124.770 -7.700 125.220 -7.590 ;
        RECT 126.170 -7.350 126.620 -7.250 ;
        RECT 128.020 -7.350 128.470 -7.250 ;
        RECT 126.170 -7.590 128.470 -7.350 ;
        RECT 126.170 -7.670 126.620 -7.590 ;
        RECT 106.680 -8.250 108.210 -8.040 ;
        RECT 108.590 -8.250 109.040 -8.160 ;
        RECT 109.420 -8.250 110.950 -8.040 ;
        RECT 120.180 -8.040 120.630 -7.760 ;
        RECT 124.000 -8.040 124.450 -7.760 ;
        RECT 127.220 -8.030 127.630 -7.590 ;
        RECT 128.020 -7.700 128.470 -7.590 ;
        RECT 129.660 -7.350 130.110 -7.250 ;
        RECT 131.510 -7.350 131.960 -7.250 ;
        RECT 129.660 -7.590 131.960 -7.350 ;
        RECT 129.660 -7.700 130.110 -7.590 ;
        RECT 130.500 -8.030 130.910 -7.590 ;
        RECT 131.510 -7.670 131.960 -7.590 ;
        RECT 132.910 -7.350 133.360 -7.280 ;
        RECT 133.960 -7.350 134.370 -6.920 ;
        RECT 134.760 -7.350 135.210 -7.250 ;
        RECT 132.910 -7.590 135.210 -7.350 ;
        RECT 132.910 -7.700 133.360 -7.590 ;
        RECT 134.760 -7.700 135.210 -7.590 ;
        RECT 136.420 -7.350 136.870 -7.250 ;
        RECT 137.260 -7.350 137.670 -6.920 ;
        RECT 140.420 -6.990 141.970 -6.770 ;
        RECT 142.350 -6.780 142.780 -6.720 ;
        RECT 143.160 -6.770 143.610 -6.720 ;
        RECT 144.210 -6.770 144.710 -6.380 ;
        RECT 143.160 -6.990 144.710 -6.770 ;
        RECT 153.920 -6.380 155.470 -6.160 ;
        RECT 153.920 -6.770 154.420 -6.380 ;
        RECT 155.020 -6.430 155.470 -6.380 ;
        RECT 155.850 -6.430 156.280 -6.370 ;
        RECT 156.660 -6.380 158.210 -6.160 ;
        RECT 160.960 -6.230 161.370 -5.800 ;
        RECT 161.760 -5.900 162.210 -5.800 ;
        RECT 163.420 -5.560 163.870 -5.450 ;
        RECT 165.270 -5.560 165.720 -5.450 ;
        RECT 163.420 -5.800 165.720 -5.560 ;
        RECT 163.420 -5.900 163.870 -5.800 ;
        RECT 164.260 -6.230 164.670 -5.800 ;
        RECT 165.270 -5.870 165.720 -5.800 ;
        RECT 166.670 -5.560 167.120 -5.480 ;
        RECT 167.720 -5.560 168.130 -5.120 ;
        RECT 168.520 -5.560 168.970 -5.450 ;
        RECT 166.670 -5.800 168.970 -5.560 ;
        RECT 166.670 -5.900 167.120 -5.800 ;
        RECT 168.520 -5.900 168.970 -5.800 ;
        RECT 170.160 -5.560 170.610 -5.450 ;
        RECT 171.000 -5.560 171.410 -5.120 ;
        RECT 174.180 -5.390 174.630 -5.110 ;
        RECT 178.000 -5.390 178.450 -5.110 ;
        RECT 187.680 -5.110 189.210 -4.900 ;
        RECT 189.590 -4.990 190.040 -4.900 ;
        RECT 190.420 -5.110 191.950 -4.900 ;
        RECT 172.010 -5.560 172.460 -5.480 ;
        RECT 170.160 -5.800 172.460 -5.560 ;
        RECT 170.160 -5.900 170.610 -5.800 ;
        RECT 172.010 -5.900 172.460 -5.800 ;
        RECT 173.410 -5.560 173.860 -5.450 ;
        RECT 175.260 -5.560 175.710 -5.450 ;
        RECT 173.410 -5.800 175.710 -5.560 ;
        RECT 173.410 -5.870 173.860 -5.800 ;
        RECT 156.660 -6.430 157.110 -6.380 ;
        RECT 155.020 -6.720 157.110 -6.430 ;
        RECT 155.020 -6.770 155.470 -6.720 ;
        RECT 138.270 -7.350 138.720 -7.280 ;
        RECT 136.420 -7.590 138.720 -7.350 ;
        RECT 136.420 -7.700 136.870 -7.590 ;
        RECT 138.270 -7.700 138.720 -7.590 ;
        RECT 139.670 -7.350 140.120 -7.250 ;
        RECT 141.520 -7.350 141.970 -7.250 ;
        RECT 139.670 -7.590 141.970 -7.350 ;
        RECT 139.670 -7.670 140.120 -7.590 ;
        RECT 120.180 -8.250 121.710 -8.040 ;
        RECT 122.090 -8.250 122.540 -8.160 ;
        RECT 122.920 -8.250 124.450 -8.040 ;
        RECT 133.680 -8.040 134.130 -7.760 ;
        RECT 137.500 -8.040 137.950 -7.760 ;
        RECT 140.720 -8.030 141.130 -7.590 ;
        RECT 141.520 -7.700 141.970 -7.590 ;
        RECT 143.160 -7.350 143.610 -7.250 ;
        RECT 145.010 -7.350 145.460 -7.250 ;
        RECT 143.160 -7.590 145.460 -7.350 ;
        RECT 143.160 -7.700 143.610 -7.590 ;
        RECT 144.000 -8.030 144.410 -7.590 ;
        RECT 145.010 -7.670 145.460 -7.590 ;
        RECT 146.410 -7.350 146.860 -7.280 ;
        RECT 147.460 -7.350 147.870 -6.920 ;
        RECT 148.260 -7.350 148.710 -7.250 ;
        RECT 146.410 -7.590 148.710 -7.350 ;
        RECT 146.410 -7.700 146.860 -7.590 ;
        RECT 148.260 -7.700 148.710 -7.590 ;
        RECT 149.920 -7.350 150.370 -7.250 ;
        RECT 150.760 -7.350 151.170 -6.920 ;
        RECT 153.920 -6.990 155.470 -6.770 ;
        RECT 155.850 -6.780 156.280 -6.720 ;
        RECT 156.660 -6.770 157.110 -6.720 ;
        RECT 157.710 -6.770 158.210 -6.380 ;
        RECT 156.660 -6.990 158.210 -6.770 ;
        RECT 167.420 -6.380 168.970 -6.160 ;
        RECT 167.420 -6.770 167.920 -6.380 ;
        RECT 168.520 -6.430 168.970 -6.380 ;
        RECT 169.350 -6.430 169.780 -6.370 ;
        RECT 170.160 -6.380 171.710 -6.160 ;
        RECT 174.460 -6.230 174.870 -5.800 ;
        RECT 175.260 -5.900 175.710 -5.800 ;
        RECT 176.920 -5.560 177.370 -5.450 ;
        RECT 178.770 -5.560 179.220 -5.450 ;
        RECT 176.920 -5.800 179.220 -5.560 ;
        RECT 176.920 -5.900 177.370 -5.800 ;
        RECT 177.760 -6.230 178.170 -5.800 ;
        RECT 178.770 -5.870 179.220 -5.800 ;
        RECT 180.170 -5.560 180.620 -5.480 ;
        RECT 181.220 -5.560 181.630 -5.120 ;
        RECT 182.020 -5.560 182.470 -5.450 ;
        RECT 180.170 -5.800 182.470 -5.560 ;
        RECT 180.170 -5.900 180.620 -5.800 ;
        RECT 182.020 -5.900 182.470 -5.800 ;
        RECT 183.660 -5.560 184.110 -5.450 ;
        RECT 184.500 -5.560 184.910 -5.120 ;
        RECT 187.680 -5.390 188.130 -5.110 ;
        RECT 191.500 -5.390 191.950 -5.110 ;
        RECT 201.180 -5.110 202.710 -4.900 ;
        RECT 203.090 -4.990 203.540 -4.900 ;
        RECT 203.920 -5.110 205.450 -4.900 ;
        RECT 185.510 -5.560 185.960 -5.480 ;
        RECT 183.660 -5.800 185.960 -5.560 ;
        RECT 183.660 -5.900 184.110 -5.800 ;
        RECT 185.510 -5.900 185.960 -5.800 ;
        RECT 186.910 -5.560 187.360 -5.450 ;
        RECT 188.760 -5.560 189.210 -5.450 ;
        RECT 186.910 -5.800 189.210 -5.560 ;
        RECT 186.910 -5.870 187.360 -5.800 ;
        RECT 170.160 -6.430 170.610 -6.380 ;
        RECT 168.520 -6.720 170.610 -6.430 ;
        RECT 168.520 -6.770 168.970 -6.720 ;
        RECT 151.770 -7.350 152.220 -7.280 ;
        RECT 149.920 -7.590 152.220 -7.350 ;
        RECT 149.920 -7.700 150.370 -7.590 ;
        RECT 151.770 -7.700 152.220 -7.590 ;
        RECT 153.170 -7.350 153.620 -7.250 ;
        RECT 155.020 -7.350 155.470 -7.250 ;
        RECT 153.170 -7.590 155.470 -7.350 ;
        RECT 153.170 -7.670 153.620 -7.590 ;
        RECT 133.680 -8.250 135.210 -8.040 ;
        RECT 135.590 -8.250 136.040 -8.160 ;
        RECT 136.420 -8.250 137.950 -8.040 ;
        RECT 147.180 -8.040 147.630 -7.760 ;
        RECT 151.000 -8.040 151.450 -7.760 ;
        RECT 154.220 -8.030 154.630 -7.590 ;
        RECT 155.020 -7.700 155.470 -7.590 ;
        RECT 156.660 -7.350 157.110 -7.250 ;
        RECT 158.510 -7.350 158.960 -7.250 ;
        RECT 156.660 -7.590 158.960 -7.350 ;
        RECT 156.660 -7.700 157.110 -7.590 ;
        RECT 157.500 -8.030 157.910 -7.590 ;
        RECT 158.510 -7.670 158.960 -7.590 ;
        RECT 159.910 -7.350 160.360 -7.280 ;
        RECT 160.960 -7.350 161.370 -6.920 ;
        RECT 161.760 -7.350 162.210 -7.250 ;
        RECT 159.910 -7.590 162.210 -7.350 ;
        RECT 159.910 -7.700 160.360 -7.590 ;
        RECT 161.760 -7.700 162.210 -7.590 ;
        RECT 163.420 -7.350 163.870 -7.250 ;
        RECT 164.260 -7.350 164.670 -6.920 ;
        RECT 167.420 -6.990 168.970 -6.770 ;
        RECT 169.350 -6.780 169.780 -6.720 ;
        RECT 170.160 -6.770 170.610 -6.720 ;
        RECT 171.210 -6.770 171.710 -6.380 ;
        RECT 170.160 -6.990 171.710 -6.770 ;
        RECT 180.920 -6.380 182.470 -6.160 ;
        RECT 180.920 -6.770 181.420 -6.380 ;
        RECT 182.020 -6.430 182.470 -6.380 ;
        RECT 182.850 -6.430 183.280 -6.370 ;
        RECT 183.660 -6.380 185.210 -6.160 ;
        RECT 187.960 -6.230 188.370 -5.800 ;
        RECT 188.760 -5.900 189.210 -5.800 ;
        RECT 190.420 -5.560 190.870 -5.450 ;
        RECT 192.270 -5.560 192.720 -5.450 ;
        RECT 190.420 -5.800 192.720 -5.560 ;
        RECT 190.420 -5.900 190.870 -5.800 ;
        RECT 191.260 -6.230 191.670 -5.800 ;
        RECT 192.270 -5.870 192.720 -5.800 ;
        RECT 193.670 -5.560 194.120 -5.480 ;
        RECT 194.720 -5.560 195.130 -5.120 ;
        RECT 195.520 -5.560 195.970 -5.450 ;
        RECT 193.670 -5.800 195.970 -5.560 ;
        RECT 193.670 -5.900 194.120 -5.800 ;
        RECT 195.520 -5.900 195.970 -5.800 ;
        RECT 197.160 -5.560 197.610 -5.450 ;
        RECT 198.000 -5.560 198.410 -5.120 ;
        RECT 201.180 -5.390 201.630 -5.110 ;
        RECT 205.000 -5.390 205.450 -5.110 ;
        RECT 214.680 -5.110 216.210 -4.900 ;
        RECT 216.590 -4.990 217.030 -4.900 ;
        RECT 199.010 -5.560 199.460 -5.480 ;
        RECT 197.160 -5.800 199.460 -5.560 ;
        RECT 197.160 -5.900 197.610 -5.800 ;
        RECT 199.010 -5.900 199.460 -5.800 ;
        RECT 200.410 -5.560 200.860 -5.450 ;
        RECT 202.260 -5.560 202.710 -5.450 ;
        RECT 200.410 -5.800 202.710 -5.560 ;
        RECT 200.410 -5.870 200.860 -5.800 ;
        RECT 183.660 -6.430 184.110 -6.380 ;
        RECT 182.020 -6.720 184.110 -6.430 ;
        RECT 182.020 -6.770 182.470 -6.720 ;
        RECT 165.270 -7.350 165.720 -7.280 ;
        RECT 163.420 -7.590 165.720 -7.350 ;
        RECT 163.420 -7.700 163.870 -7.590 ;
        RECT 165.270 -7.700 165.720 -7.590 ;
        RECT 166.670 -7.350 167.120 -7.250 ;
        RECT 168.520 -7.350 168.970 -7.250 ;
        RECT 166.670 -7.590 168.970 -7.350 ;
        RECT 166.670 -7.670 167.120 -7.590 ;
        RECT 147.180 -8.250 148.710 -8.040 ;
        RECT 149.090 -8.250 149.540 -8.160 ;
        RECT 149.920 -8.250 151.450 -8.040 ;
        RECT 160.680 -8.040 161.130 -7.760 ;
        RECT 164.500 -8.040 164.950 -7.760 ;
        RECT 167.720 -8.030 168.130 -7.590 ;
        RECT 168.520 -7.700 168.970 -7.590 ;
        RECT 170.160 -7.350 170.610 -7.250 ;
        RECT 172.010 -7.350 172.460 -7.250 ;
        RECT 170.160 -7.590 172.460 -7.350 ;
        RECT 170.160 -7.700 170.610 -7.590 ;
        RECT 171.000 -8.030 171.410 -7.590 ;
        RECT 172.010 -7.670 172.460 -7.590 ;
        RECT 173.410 -7.350 173.860 -7.280 ;
        RECT 174.460 -7.350 174.870 -6.920 ;
        RECT 175.260 -7.350 175.710 -7.250 ;
        RECT 173.410 -7.590 175.710 -7.350 ;
        RECT 173.410 -7.700 173.860 -7.590 ;
        RECT 175.260 -7.700 175.710 -7.590 ;
        RECT 176.920 -7.350 177.370 -7.250 ;
        RECT 177.760 -7.350 178.170 -6.920 ;
        RECT 180.920 -6.990 182.470 -6.770 ;
        RECT 182.850 -6.780 183.280 -6.720 ;
        RECT 183.660 -6.770 184.110 -6.720 ;
        RECT 184.710 -6.770 185.210 -6.380 ;
        RECT 183.660 -6.990 185.210 -6.770 ;
        RECT 194.420 -6.380 195.970 -6.160 ;
        RECT 194.420 -6.770 194.920 -6.380 ;
        RECT 195.520 -6.430 195.970 -6.380 ;
        RECT 196.350 -6.430 196.780 -6.370 ;
        RECT 197.160 -6.380 198.710 -6.160 ;
        RECT 201.460 -6.230 201.870 -5.800 ;
        RECT 202.260 -5.900 202.710 -5.800 ;
        RECT 203.920 -5.560 204.370 -5.450 ;
        RECT 205.770 -5.560 206.220 -5.450 ;
        RECT 203.920 -5.800 206.220 -5.560 ;
        RECT 203.920 -5.900 204.370 -5.800 ;
        RECT 204.760 -6.230 205.170 -5.800 ;
        RECT 205.770 -5.870 206.220 -5.800 ;
        RECT 207.170 -5.560 207.620 -5.480 ;
        RECT 208.220 -5.560 208.630 -5.120 ;
        RECT 209.020 -5.560 209.470 -5.450 ;
        RECT 207.170 -5.800 209.470 -5.560 ;
        RECT 207.170 -5.900 207.620 -5.800 ;
        RECT 209.020 -5.900 209.470 -5.800 ;
        RECT 210.660 -5.560 211.110 -5.450 ;
        RECT 211.500 -5.560 211.910 -5.120 ;
        RECT 214.680 -5.390 215.130 -5.110 ;
        RECT 212.510 -5.560 212.960 -5.480 ;
        RECT 210.660 -5.800 212.960 -5.560 ;
        RECT 210.660 -5.900 211.110 -5.800 ;
        RECT 212.510 -5.900 212.960 -5.800 ;
        RECT 213.910 -5.560 214.360 -5.450 ;
        RECT 215.760 -5.560 216.210 -5.450 ;
        RECT 213.910 -5.800 216.210 -5.560 ;
        RECT 213.910 -5.870 214.360 -5.800 ;
        RECT 197.160 -6.430 197.610 -6.380 ;
        RECT 195.520 -6.720 197.610 -6.430 ;
        RECT 195.520 -6.770 195.970 -6.720 ;
        RECT 178.770 -7.350 179.220 -7.280 ;
        RECT 176.920 -7.590 179.220 -7.350 ;
        RECT 176.920 -7.700 177.370 -7.590 ;
        RECT 178.770 -7.700 179.220 -7.590 ;
        RECT 180.170 -7.350 180.620 -7.250 ;
        RECT 182.020 -7.350 182.470 -7.250 ;
        RECT 180.170 -7.590 182.470 -7.350 ;
        RECT 180.170 -7.670 180.620 -7.590 ;
        RECT 160.680 -8.250 162.210 -8.040 ;
        RECT 162.590 -8.250 163.040 -8.160 ;
        RECT 163.420 -8.250 164.950 -8.040 ;
        RECT 174.180 -8.040 174.630 -7.760 ;
        RECT 178.000 -8.040 178.450 -7.760 ;
        RECT 181.220 -8.030 181.630 -7.590 ;
        RECT 182.020 -7.700 182.470 -7.590 ;
        RECT 183.660 -7.350 184.110 -7.250 ;
        RECT 185.510 -7.350 185.960 -7.250 ;
        RECT 183.660 -7.590 185.960 -7.350 ;
        RECT 183.660 -7.700 184.110 -7.590 ;
        RECT 184.500 -8.030 184.910 -7.590 ;
        RECT 185.510 -7.670 185.960 -7.590 ;
        RECT 186.910 -7.350 187.360 -7.280 ;
        RECT 187.960 -7.350 188.370 -6.920 ;
        RECT 188.760 -7.350 189.210 -7.250 ;
        RECT 186.910 -7.590 189.210 -7.350 ;
        RECT 186.910 -7.700 187.360 -7.590 ;
        RECT 188.760 -7.700 189.210 -7.590 ;
        RECT 190.420 -7.350 190.870 -7.250 ;
        RECT 191.260 -7.350 191.670 -6.920 ;
        RECT 194.420 -6.990 195.970 -6.770 ;
        RECT 196.350 -6.780 196.780 -6.720 ;
        RECT 197.160 -6.770 197.610 -6.720 ;
        RECT 198.210 -6.770 198.710 -6.380 ;
        RECT 197.160 -6.990 198.710 -6.770 ;
        RECT 207.920 -6.380 209.470 -6.160 ;
        RECT 207.920 -6.770 208.420 -6.380 ;
        RECT 209.020 -6.430 209.470 -6.380 ;
        RECT 209.850 -6.430 210.280 -6.370 ;
        RECT 210.660 -6.380 212.210 -6.160 ;
        RECT 214.960 -6.230 215.370 -5.800 ;
        RECT 215.760 -5.900 216.210 -5.800 ;
        RECT 210.660 -6.430 211.110 -6.380 ;
        RECT 209.020 -6.720 211.110 -6.430 ;
        RECT 209.020 -6.770 209.470 -6.720 ;
        RECT 192.270 -7.350 192.720 -7.280 ;
        RECT 190.420 -7.590 192.720 -7.350 ;
        RECT 190.420 -7.700 190.870 -7.590 ;
        RECT 192.270 -7.700 192.720 -7.590 ;
        RECT 193.670 -7.350 194.120 -7.250 ;
        RECT 195.520 -7.350 195.970 -7.250 ;
        RECT 193.670 -7.590 195.970 -7.350 ;
        RECT 193.670 -7.670 194.120 -7.590 ;
        RECT 174.180 -8.250 175.710 -8.040 ;
        RECT 176.090 -8.250 176.540 -8.160 ;
        RECT 176.920 -8.250 178.450 -8.040 ;
        RECT 187.680 -8.040 188.130 -7.760 ;
        RECT 191.500 -8.040 191.950 -7.760 ;
        RECT 194.720 -8.030 195.130 -7.590 ;
        RECT 195.520 -7.700 195.970 -7.590 ;
        RECT 197.160 -7.350 197.610 -7.250 ;
        RECT 199.010 -7.350 199.460 -7.250 ;
        RECT 197.160 -7.590 199.460 -7.350 ;
        RECT 197.160 -7.700 197.610 -7.590 ;
        RECT 198.000 -8.030 198.410 -7.590 ;
        RECT 199.010 -7.670 199.460 -7.590 ;
        RECT 200.410 -7.350 200.860 -7.280 ;
        RECT 201.460 -7.350 201.870 -6.920 ;
        RECT 202.260 -7.350 202.710 -7.250 ;
        RECT 200.410 -7.590 202.710 -7.350 ;
        RECT 200.410 -7.700 200.860 -7.590 ;
        RECT 202.260 -7.700 202.710 -7.590 ;
        RECT 203.920 -7.350 204.370 -7.250 ;
        RECT 204.760 -7.350 205.170 -6.920 ;
        RECT 207.920 -6.990 209.470 -6.770 ;
        RECT 209.850 -6.780 210.280 -6.720 ;
        RECT 210.660 -6.770 211.110 -6.720 ;
        RECT 211.710 -6.770 212.210 -6.380 ;
        RECT 210.660 -6.990 212.210 -6.770 ;
        RECT 205.770 -7.350 206.220 -7.280 ;
        RECT 203.920 -7.590 206.220 -7.350 ;
        RECT 203.920 -7.700 204.370 -7.590 ;
        RECT 205.770 -7.700 206.220 -7.590 ;
        RECT 207.170 -7.350 207.620 -7.250 ;
        RECT 209.020 -7.350 209.470 -7.250 ;
        RECT 207.170 -7.590 209.470 -7.350 ;
        RECT 207.170 -7.670 207.620 -7.590 ;
        RECT 187.680 -8.250 189.210 -8.040 ;
        RECT 189.590 -8.250 190.040 -8.160 ;
        RECT 190.420 -8.250 191.950 -8.040 ;
        RECT 201.180 -8.040 201.630 -7.760 ;
        RECT 205.000 -8.040 205.450 -7.760 ;
        RECT 208.220 -8.030 208.630 -7.590 ;
        RECT 209.020 -7.700 209.470 -7.590 ;
        RECT 210.660 -7.350 211.110 -7.250 ;
        RECT 212.510 -7.350 212.960 -7.250 ;
        RECT 210.660 -7.590 212.960 -7.350 ;
        RECT 210.660 -7.700 211.110 -7.590 ;
        RECT 211.500 -8.030 211.910 -7.590 ;
        RECT 212.510 -7.670 212.960 -7.590 ;
        RECT 213.910 -7.350 214.360 -7.280 ;
        RECT 214.960 -7.350 215.370 -6.920 ;
        RECT 215.760 -7.350 216.210 -7.250 ;
        RECT 213.910 -7.590 216.210 -7.350 ;
        RECT 213.910 -7.700 214.360 -7.590 ;
        RECT 215.760 -7.700 216.210 -7.590 ;
        RECT 201.180 -8.250 202.710 -8.040 ;
        RECT 203.090 -8.250 203.540 -8.160 ;
        RECT 203.920 -8.250 205.450 -8.040 ;
        RECT 214.680 -8.040 215.130 -7.760 ;
        RECT 214.680 -8.250 216.210 -8.040 ;
        RECT 216.590 -8.250 217.030 -8.160 ;
        RECT 13.260 -8.510 15.370 -8.250 ;
        RECT 26.760 -8.510 28.870 -8.250 ;
        RECT 40.260 -8.510 42.370 -8.250 ;
        RECT 53.760 -8.510 55.870 -8.250 ;
        RECT 67.260 -8.510 69.370 -8.250 ;
        RECT 80.760 -8.510 82.870 -8.250 ;
        RECT 94.260 -8.510 96.370 -8.250 ;
        RECT 107.760 -8.510 109.870 -8.250 ;
        RECT 121.260 -8.510 123.370 -8.250 ;
        RECT 134.760 -8.510 136.870 -8.250 ;
        RECT 148.260 -8.510 150.370 -8.250 ;
        RECT 161.760 -8.510 163.870 -8.250 ;
        RECT 175.260 -8.510 177.370 -8.250 ;
        RECT 188.760 -8.510 190.870 -8.250 ;
        RECT 202.260 -8.510 204.370 -8.250 ;
        RECT 215.760 -8.310 217.030 -8.250 ;
        RECT 215.760 -8.500 217.240 -8.310 ;
        RECT 215.760 -8.510 217.030 -8.500 ;
        RECT 12.180 -8.720 13.710 -8.510 ;
        RECT 14.090 -8.600 14.540 -8.510 ;
        RECT 14.920 -8.720 16.450 -8.510 ;
        RECT 1.420 -9.170 1.870 -9.060 ;
        RECT 3.270 -9.170 3.720 -9.060 ;
        RECT 1.420 -9.410 3.720 -9.170 ;
        RECT 1.420 -9.510 1.870 -9.410 ;
        RECT 2.260 -9.840 2.670 -9.410 ;
        RECT 3.270 -9.480 3.720 -9.410 ;
        RECT 4.670 -9.170 5.120 -9.090 ;
        RECT 5.720 -9.170 6.130 -8.730 ;
        RECT 6.520 -9.170 6.970 -9.060 ;
        RECT 4.670 -9.410 6.970 -9.170 ;
        RECT 4.670 -9.510 5.120 -9.410 ;
        RECT 6.520 -9.510 6.970 -9.410 ;
        RECT 8.160 -9.170 8.610 -9.060 ;
        RECT 9.000 -9.170 9.410 -8.730 ;
        RECT 12.180 -9.000 12.630 -8.720 ;
        RECT 16.000 -9.000 16.450 -8.720 ;
        RECT 25.680 -8.720 27.210 -8.510 ;
        RECT 27.590 -8.600 28.040 -8.510 ;
        RECT 28.420 -8.720 29.950 -8.510 ;
        RECT 10.010 -9.170 10.460 -9.090 ;
        RECT 8.160 -9.410 10.460 -9.170 ;
        RECT 8.160 -9.510 8.610 -9.410 ;
        RECT 10.010 -9.510 10.460 -9.410 ;
        RECT 11.410 -9.170 11.860 -9.060 ;
        RECT 13.260 -9.170 13.710 -9.060 ;
        RECT 11.410 -9.410 13.710 -9.170 ;
        RECT 11.410 -9.480 11.860 -9.410 ;
        RECT 5.420 -9.990 6.970 -9.770 ;
        RECT 5.420 -10.380 5.920 -9.990 ;
        RECT 6.520 -10.040 6.970 -9.990 ;
        RECT 7.350 -10.040 7.780 -9.980 ;
        RECT 8.160 -9.990 9.710 -9.770 ;
        RECT 12.460 -9.840 12.870 -9.410 ;
        RECT 13.260 -9.510 13.710 -9.410 ;
        RECT 14.920 -9.170 15.370 -9.060 ;
        RECT 16.770 -9.170 17.220 -9.060 ;
        RECT 14.920 -9.410 17.220 -9.170 ;
        RECT 14.920 -9.510 15.370 -9.410 ;
        RECT 15.760 -9.840 16.170 -9.410 ;
        RECT 16.770 -9.480 17.220 -9.410 ;
        RECT 18.170 -9.170 18.620 -9.090 ;
        RECT 19.220 -9.170 19.630 -8.730 ;
        RECT 20.020 -9.170 20.470 -9.060 ;
        RECT 18.170 -9.410 20.470 -9.170 ;
        RECT 18.170 -9.510 18.620 -9.410 ;
        RECT 20.020 -9.510 20.470 -9.410 ;
        RECT 21.660 -9.170 22.110 -9.060 ;
        RECT 22.500 -9.170 22.910 -8.730 ;
        RECT 25.680 -9.000 26.130 -8.720 ;
        RECT 29.500 -9.000 29.950 -8.720 ;
        RECT 39.180 -8.720 40.710 -8.510 ;
        RECT 41.090 -8.600 41.540 -8.510 ;
        RECT 41.920 -8.720 43.450 -8.510 ;
        RECT 23.510 -9.170 23.960 -9.090 ;
        RECT 21.660 -9.410 23.960 -9.170 ;
        RECT 21.660 -9.510 22.110 -9.410 ;
        RECT 23.510 -9.510 23.960 -9.410 ;
        RECT 24.910 -9.170 25.360 -9.060 ;
        RECT 26.760 -9.170 27.210 -9.060 ;
        RECT 24.910 -9.410 27.210 -9.170 ;
        RECT 24.910 -9.480 25.360 -9.410 ;
        RECT 8.160 -10.040 8.610 -9.990 ;
        RECT 6.520 -10.330 8.610 -10.040 ;
        RECT 6.520 -10.380 6.970 -10.330 ;
        RECT 1.420 -10.960 1.870 -10.860 ;
        RECT 2.260 -10.960 2.670 -10.530 ;
        RECT 5.420 -10.600 6.970 -10.380 ;
        RECT 7.350 -10.390 7.780 -10.330 ;
        RECT 8.160 -10.380 8.610 -10.330 ;
        RECT 9.210 -10.380 9.710 -9.990 ;
        RECT 8.160 -10.600 9.710 -10.380 ;
        RECT 18.920 -9.990 20.470 -9.770 ;
        RECT 18.920 -10.380 19.420 -9.990 ;
        RECT 20.020 -10.040 20.470 -9.990 ;
        RECT 20.850 -10.040 21.280 -9.980 ;
        RECT 21.660 -9.990 23.210 -9.770 ;
        RECT 25.960 -9.840 26.370 -9.410 ;
        RECT 26.760 -9.510 27.210 -9.410 ;
        RECT 28.420 -9.170 28.870 -9.060 ;
        RECT 30.270 -9.170 30.720 -9.060 ;
        RECT 28.420 -9.410 30.720 -9.170 ;
        RECT 28.420 -9.510 28.870 -9.410 ;
        RECT 29.260 -9.840 29.670 -9.410 ;
        RECT 30.270 -9.480 30.720 -9.410 ;
        RECT 31.670 -9.170 32.120 -9.090 ;
        RECT 32.720 -9.170 33.130 -8.730 ;
        RECT 33.520 -9.170 33.970 -9.060 ;
        RECT 31.670 -9.410 33.970 -9.170 ;
        RECT 31.670 -9.510 32.120 -9.410 ;
        RECT 33.520 -9.510 33.970 -9.410 ;
        RECT 35.160 -9.170 35.610 -9.060 ;
        RECT 36.000 -9.170 36.410 -8.730 ;
        RECT 39.180 -9.000 39.630 -8.720 ;
        RECT 43.000 -9.000 43.450 -8.720 ;
        RECT 52.680 -8.720 54.210 -8.510 ;
        RECT 54.590 -8.600 55.040 -8.510 ;
        RECT 55.420 -8.720 56.950 -8.510 ;
        RECT 37.010 -9.170 37.460 -9.090 ;
        RECT 35.160 -9.410 37.460 -9.170 ;
        RECT 35.160 -9.510 35.610 -9.410 ;
        RECT 37.010 -9.510 37.460 -9.410 ;
        RECT 38.410 -9.170 38.860 -9.060 ;
        RECT 40.260 -9.170 40.710 -9.060 ;
        RECT 38.410 -9.410 40.710 -9.170 ;
        RECT 38.410 -9.480 38.860 -9.410 ;
        RECT 21.660 -10.040 22.110 -9.990 ;
        RECT 20.020 -10.330 22.110 -10.040 ;
        RECT 20.020 -10.380 20.470 -10.330 ;
        RECT 3.270 -10.960 3.720 -10.890 ;
        RECT 1.420 -11.200 3.720 -10.960 ;
        RECT 1.420 -11.310 1.870 -11.200 ;
        RECT 3.270 -11.310 3.720 -11.200 ;
        RECT 4.670 -10.960 5.120 -10.860 ;
        RECT 6.520 -10.960 6.970 -10.860 ;
        RECT 4.670 -11.200 6.970 -10.960 ;
        RECT 4.670 -11.280 5.120 -11.200 ;
        RECT 5.720 -11.640 6.130 -11.200 ;
        RECT 6.520 -11.310 6.970 -11.200 ;
        RECT 8.160 -10.960 8.610 -10.860 ;
        RECT 10.010 -10.960 10.460 -10.860 ;
        RECT 8.160 -11.200 10.460 -10.960 ;
        RECT 8.160 -11.310 8.610 -11.200 ;
        RECT 9.000 -11.640 9.410 -11.200 ;
        RECT 10.010 -11.280 10.460 -11.200 ;
        RECT 11.410 -10.960 11.860 -10.890 ;
        RECT 12.460 -10.960 12.870 -10.530 ;
        RECT 13.260 -10.960 13.710 -10.860 ;
        RECT 11.410 -11.200 13.710 -10.960 ;
        RECT 11.410 -11.310 11.860 -11.200 ;
        RECT 13.260 -11.310 13.710 -11.200 ;
        RECT 14.920 -10.960 15.370 -10.860 ;
        RECT 15.760 -10.960 16.170 -10.530 ;
        RECT 18.920 -10.600 20.470 -10.380 ;
        RECT 20.850 -10.390 21.280 -10.330 ;
        RECT 21.660 -10.380 22.110 -10.330 ;
        RECT 22.710 -10.380 23.210 -9.990 ;
        RECT 21.660 -10.600 23.210 -10.380 ;
        RECT 32.420 -9.990 33.970 -9.770 ;
        RECT 32.420 -10.380 32.920 -9.990 ;
        RECT 33.520 -10.040 33.970 -9.990 ;
        RECT 34.350 -10.040 34.780 -9.980 ;
        RECT 35.160 -9.990 36.710 -9.770 ;
        RECT 39.460 -9.840 39.870 -9.410 ;
        RECT 40.260 -9.510 40.710 -9.410 ;
        RECT 41.920 -9.170 42.370 -9.060 ;
        RECT 43.770 -9.170 44.220 -9.060 ;
        RECT 41.920 -9.410 44.220 -9.170 ;
        RECT 41.920 -9.510 42.370 -9.410 ;
        RECT 42.760 -9.840 43.170 -9.410 ;
        RECT 43.770 -9.480 44.220 -9.410 ;
        RECT 45.170 -9.170 45.620 -9.090 ;
        RECT 46.220 -9.170 46.630 -8.730 ;
        RECT 47.020 -9.170 47.470 -9.060 ;
        RECT 45.170 -9.410 47.470 -9.170 ;
        RECT 45.170 -9.510 45.620 -9.410 ;
        RECT 47.020 -9.510 47.470 -9.410 ;
        RECT 48.660 -9.170 49.110 -9.060 ;
        RECT 49.500 -9.170 49.910 -8.730 ;
        RECT 52.680 -9.000 53.130 -8.720 ;
        RECT 56.500 -9.000 56.950 -8.720 ;
        RECT 66.180 -8.720 67.710 -8.510 ;
        RECT 68.090 -8.600 68.540 -8.510 ;
        RECT 68.920 -8.720 70.450 -8.510 ;
        RECT 50.510 -9.170 50.960 -9.090 ;
        RECT 48.660 -9.410 50.960 -9.170 ;
        RECT 48.660 -9.510 49.110 -9.410 ;
        RECT 50.510 -9.510 50.960 -9.410 ;
        RECT 51.910 -9.170 52.360 -9.060 ;
        RECT 53.760 -9.170 54.210 -9.060 ;
        RECT 51.910 -9.410 54.210 -9.170 ;
        RECT 51.910 -9.480 52.360 -9.410 ;
        RECT 35.160 -10.040 35.610 -9.990 ;
        RECT 33.520 -10.330 35.610 -10.040 ;
        RECT 33.520 -10.380 33.970 -10.330 ;
        RECT 16.770 -10.960 17.220 -10.890 ;
        RECT 14.920 -11.200 17.220 -10.960 ;
        RECT 14.920 -11.310 15.370 -11.200 ;
        RECT 16.770 -11.310 17.220 -11.200 ;
        RECT 18.170 -10.960 18.620 -10.860 ;
        RECT 20.020 -10.960 20.470 -10.860 ;
        RECT 18.170 -11.200 20.470 -10.960 ;
        RECT 18.170 -11.280 18.620 -11.200 ;
        RECT 12.180 -11.650 12.630 -11.370 ;
        RECT 16.000 -11.650 16.450 -11.370 ;
        RECT 19.220 -11.640 19.630 -11.200 ;
        RECT 20.020 -11.310 20.470 -11.200 ;
        RECT 21.660 -10.960 22.110 -10.860 ;
        RECT 23.510 -10.960 23.960 -10.860 ;
        RECT 21.660 -11.200 23.960 -10.960 ;
        RECT 21.660 -11.310 22.110 -11.200 ;
        RECT 22.500 -11.640 22.910 -11.200 ;
        RECT 23.510 -11.280 23.960 -11.200 ;
        RECT 24.910 -10.960 25.360 -10.890 ;
        RECT 25.960 -10.960 26.370 -10.530 ;
        RECT 26.760 -10.960 27.210 -10.860 ;
        RECT 24.910 -11.200 27.210 -10.960 ;
        RECT 24.910 -11.310 25.360 -11.200 ;
        RECT 26.760 -11.310 27.210 -11.200 ;
        RECT 28.420 -10.960 28.870 -10.860 ;
        RECT 29.260 -10.960 29.670 -10.530 ;
        RECT 32.420 -10.600 33.970 -10.380 ;
        RECT 34.350 -10.390 34.780 -10.330 ;
        RECT 35.160 -10.380 35.610 -10.330 ;
        RECT 36.210 -10.380 36.710 -9.990 ;
        RECT 35.160 -10.600 36.710 -10.380 ;
        RECT 45.920 -9.990 47.470 -9.770 ;
        RECT 45.920 -10.380 46.420 -9.990 ;
        RECT 47.020 -10.040 47.470 -9.990 ;
        RECT 47.850 -10.040 48.280 -9.980 ;
        RECT 48.660 -9.990 50.210 -9.770 ;
        RECT 52.960 -9.840 53.370 -9.410 ;
        RECT 53.760 -9.510 54.210 -9.410 ;
        RECT 55.420 -9.170 55.870 -9.060 ;
        RECT 57.270 -9.170 57.720 -9.060 ;
        RECT 55.420 -9.410 57.720 -9.170 ;
        RECT 55.420 -9.510 55.870 -9.410 ;
        RECT 56.260 -9.840 56.670 -9.410 ;
        RECT 57.270 -9.480 57.720 -9.410 ;
        RECT 58.670 -9.170 59.120 -9.090 ;
        RECT 59.720 -9.170 60.130 -8.730 ;
        RECT 60.520 -9.170 60.970 -9.060 ;
        RECT 58.670 -9.410 60.970 -9.170 ;
        RECT 58.670 -9.510 59.120 -9.410 ;
        RECT 60.520 -9.510 60.970 -9.410 ;
        RECT 62.160 -9.170 62.610 -9.060 ;
        RECT 63.000 -9.170 63.410 -8.730 ;
        RECT 66.180 -9.000 66.630 -8.720 ;
        RECT 70.000 -9.000 70.450 -8.720 ;
        RECT 79.680 -8.720 81.210 -8.510 ;
        RECT 81.590 -8.600 82.040 -8.510 ;
        RECT 82.420 -8.720 83.950 -8.510 ;
        RECT 64.010 -9.170 64.460 -9.090 ;
        RECT 62.160 -9.410 64.460 -9.170 ;
        RECT 62.160 -9.510 62.610 -9.410 ;
        RECT 64.010 -9.510 64.460 -9.410 ;
        RECT 65.410 -9.170 65.860 -9.060 ;
        RECT 67.260 -9.170 67.710 -9.060 ;
        RECT 65.410 -9.410 67.710 -9.170 ;
        RECT 65.410 -9.480 65.860 -9.410 ;
        RECT 48.660 -10.040 49.110 -9.990 ;
        RECT 47.020 -10.330 49.110 -10.040 ;
        RECT 47.020 -10.380 47.470 -10.330 ;
        RECT 30.270 -10.960 30.720 -10.890 ;
        RECT 28.420 -11.200 30.720 -10.960 ;
        RECT 28.420 -11.310 28.870 -11.200 ;
        RECT 30.270 -11.310 30.720 -11.200 ;
        RECT 31.670 -10.960 32.120 -10.860 ;
        RECT 33.520 -10.960 33.970 -10.860 ;
        RECT 31.670 -11.200 33.970 -10.960 ;
        RECT 31.670 -11.280 32.120 -11.200 ;
        RECT 12.180 -11.860 13.710 -11.650 ;
        RECT 14.090 -11.860 14.540 -11.770 ;
        RECT 14.920 -11.860 16.450 -11.650 ;
        RECT 25.680 -11.650 26.130 -11.370 ;
        RECT 29.500 -11.650 29.950 -11.370 ;
        RECT 32.720 -11.640 33.130 -11.200 ;
        RECT 33.520 -11.310 33.970 -11.200 ;
        RECT 35.160 -10.960 35.610 -10.860 ;
        RECT 37.010 -10.960 37.460 -10.860 ;
        RECT 35.160 -11.200 37.460 -10.960 ;
        RECT 35.160 -11.310 35.610 -11.200 ;
        RECT 36.000 -11.640 36.410 -11.200 ;
        RECT 37.010 -11.280 37.460 -11.200 ;
        RECT 38.410 -10.960 38.860 -10.890 ;
        RECT 39.460 -10.960 39.870 -10.530 ;
        RECT 40.260 -10.960 40.710 -10.860 ;
        RECT 38.410 -11.200 40.710 -10.960 ;
        RECT 38.410 -11.310 38.860 -11.200 ;
        RECT 40.260 -11.310 40.710 -11.200 ;
        RECT 41.920 -10.960 42.370 -10.860 ;
        RECT 42.760 -10.960 43.170 -10.530 ;
        RECT 45.920 -10.600 47.470 -10.380 ;
        RECT 47.850 -10.390 48.280 -10.330 ;
        RECT 48.660 -10.380 49.110 -10.330 ;
        RECT 49.710 -10.380 50.210 -9.990 ;
        RECT 48.660 -10.600 50.210 -10.380 ;
        RECT 59.420 -9.990 60.970 -9.770 ;
        RECT 59.420 -10.380 59.920 -9.990 ;
        RECT 60.520 -10.040 60.970 -9.990 ;
        RECT 61.350 -10.040 61.780 -9.980 ;
        RECT 62.160 -9.990 63.710 -9.770 ;
        RECT 66.460 -9.840 66.870 -9.410 ;
        RECT 67.260 -9.510 67.710 -9.410 ;
        RECT 68.920 -9.170 69.370 -9.060 ;
        RECT 70.770 -9.170 71.220 -9.060 ;
        RECT 68.920 -9.410 71.220 -9.170 ;
        RECT 68.920 -9.510 69.370 -9.410 ;
        RECT 69.760 -9.840 70.170 -9.410 ;
        RECT 70.770 -9.480 71.220 -9.410 ;
        RECT 72.170 -9.170 72.620 -9.090 ;
        RECT 73.220 -9.170 73.630 -8.730 ;
        RECT 74.020 -9.170 74.470 -9.060 ;
        RECT 72.170 -9.410 74.470 -9.170 ;
        RECT 72.170 -9.510 72.620 -9.410 ;
        RECT 74.020 -9.510 74.470 -9.410 ;
        RECT 75.660 -9.170 76.110 -9.060 ;
        RECT 76.500 -9.170 76.910 -8.730 ;
        RECT 79.680 -9.000 80.130 -8.720 ;
        RECT 83.500 -9.000 83.950 -8.720 ;
        RECT 93.180 -8.720 94.710 -8.510 ;
        RECT 95.090 -8.600 95.540 -8.510 ;
        RECT 95.920 -8.720 97.450 -8.510 ;
        RECT 77.510 -9.170 77.960 -9.090 ;
        RECT 75.660 -9.410 77.960 -9.170 ;
        RECT 75.660 -9.510 76.110 -9.410 ;
        RECT 77.510 -9.510 77.960 -9.410 ;
        RECT 78.910 -9.170 79.360 -9.060 ;
        RECT 80.760 -9.170 81.210 -9.060 ;
        RECT 78.910 -9.410 81.210 -9.170 ;
        RECT 78.910 -9.480 79.360 -9.410 ;
        RECT 62.160 -10.040 62.610 -9.990 ;
        RECT 60.520 -10.330 62.610 -10.040 ;
        RECT 60.520 -10.380 60.970 -10.330 ;
        RECT 43.770 -10.960 44.220 -10.890 ;
        RECT 41.920 -11.200 44.220 -10.960 ;
        RECT 41.920 -11.310 42.370 -11.200 ;
        RECT 43.770 -11.310 44.220 -11.200 ;
        RECT 45.170 -10.960 45.620 -10.860 ;
        RECT 47.020 -10.960 47.470 -10.860 ;
        RECT 45.170 -11.200 47.470 -10.960 ;
        RECT 45.170 -11.280 45.620 -11.200 ;
        RECT 25.680 -11.860 27.210 -11.650 ;
        RECT 27.590 -11.860 28.040 -11.770 ;
        RECT 28.420 -11.860 29.950 -11.650 ;
        RECT 39.180 -11.650 39.630 -11.370 ;
        RECT 43.000 -11.650 43.450 -11.370 ;
        RECT 46.220 -11.640 46.630 -11.200 ;
        RECT 47.020 -11.310 47.470 -11.200 ;
        RECT 48.660 -10.960 49.110 -10.860 ;
        RECT 50.510 -10.960 50.960 -10.860 ;
        RECT 48.660 -11.200 50.960 -10.960 ;
        RECT 48.660 -11.310 49.110 -11.200 ;
        RECT 49.500 -11.640 49.910 -11.200 ;
        RECT 50.510 -11.280 50.960 -11.200 ;
        RECT 51.910 -10.960 52.360 -10.890 ;
        RECT 52.960 -10.960 53.370 -10.530 ;
        RECT 53.760 -10.960 54.210 -10.860 ;
        RECT 51.910 -11.200 54.210 -10.960 ;
        RECT 51.910 -11.310 52.360 -11.200 ;
        RECT 53.760 -11.310 54.210 -11.200 ;
        RECT 55.420 -10.960 55.870 -10.860 ;
        RECT 56.260 -10.960 56.670 -10.530 ;
        RECT 59.420 -10.600 60.970 -10.380 ;
        RECT 61.350 -10.390 61.780 -10.330 ;
        RECT 62.160 -10.380 62.610 -10.330 ;
        RECT 63.210 -10.380 63.710 -9.990 ;
        RECT 62.160 -10.600 63.710 -10.380 ;
        RECT 72.920 -9.990 74.470 -9.770 ;
        RECT 72.920 -10.380 73.420 -9.990 ;
        RECT 74.020 -10.040 74.470 -9.990 ;
        RECT 74.850 -10.040 75.280 -9.980 ;
        RECT 75.660 -9.990 77.210 -9.770 ;
        RECT 79.960 -9.840 80.370 -9.410 ;
        RECT 80.760 -9.510 81.210 -9.410 ;
        RECT 82.420 -9.170 82.870 -9.060 ;
        RECT 84.270 -9.170 84.720 -9.060 ;
        RECT 82.420 -9.410 84.720 -9.170 ;
        RECT 82.420 -9.510 82.870 -9.410 ;
        RECT 83.260 -9.840 83.670 -9.410 ;
        RECT 84.270 -9.480 84.720 -9.410 ;
        RECT 85.670 -9.170 86.120 -9.090 ;
        RECT 86.720 -9.170 87.130 -8.730 ;
        RECT 87.520 -9.170 87.970 -9.060 ;
        RECT 85.670 -9.410 87.970 -9.170 ;
        RECT 85.670 -9.510 86.120 -9.410 ;
        RECT 87.520 -9.510 87.970 -9.410 ;
        RECT 89.160 -9.170 89.610 -9.060 ;
        RECT 90.000 -9.170 90.410 -8.730 ;
        RECT 93.180 -9.000 93.630 -8.720 ;
        RECT 97.000 -9.000 97.450 -8.720 ;
        RECT 106.680 -8.720 108.210 -8.510 ;
        RECT 108.590 -8.600 109.040 -8.510 ;
        RECT 109.420 -8.720 110.950 -8.510 ;
        RECT 91.010 -9.170 91.460 -9.090 ;
        RECT 89.160 -9.410 91.460 -9.170 ;
        RECT 89.160 -9.510 89.610 -9.410 ;
        RECT 91.010 -9.510 91.460 -9.410 ;
        RECT 92.410 -9.170 92.860 -9.060 ;
        RECT 94.260 -9.170 94.710 -9.060 ;
        RECT 92.410 -9.410 94.710 -9.170 ;
        RECT 92.410 -9.480 92.860 -9.410 ;
        RECT 75.660 -10.040 76.110 -9.990 ;
        RECT 74.020 -10.330 76.110 -10.040 ;
        RECT 74.020 -10.380 74.470 -10.330 ;
        RECT 57.270 -10.960 57.720 -10.890 ;
        RECT 55.420 -11.200 57.720 -10.960 ;
        RECT 55.420 -11.310 55.870 -11.200 ;
        RECT 57.270 -11.310 57.720 -11.200 ;
        RECT 58.670 -10.960 59.120 -10.860 ;
        RECT 60.520 -10.960 60.970 -10.860 ;
        RECT 58.670 -11.200 60.970 -10.960 ;
        RECT 58.670 -11.280 59.120 -11.200 ;
        RECT 39.180 -11.860 40.710 -11.650 ;
        RECT 41.090 -11.860 41.540 -11.770 ;
        RECT 41.920 -11.860 43.450 -11.650 ;
        RECT 52.680 -11.650 53.130 -11.370 ;
        RECT 56.500 -11.650 56.950 -11.370 ;
        RECT 59.720 -11.640 60.130 -11.200 ;
        RECT 60.520 -11.310 60.970 -11.200 ;
        RECT 62.160 -10.960 62.610 -10.860 ;
        RECT 64.010 -10.960 64.460 -10.860 ;
        RECT 62.160 -11.200 64.460 -10.960 ;
        RECT 62.160 -11.310 62.610 -11.200 ;
        RECT 63.000 -11.640 63.410 -11.200 ;
        RECT 64.010 -11.280 64.460 -11.200 ;
        RECT 65.410 -10.960 65.860 -10.890 ;
        RECT 66.460 -10.960 66.870 -10.530 ;
        RECT 67.260 -10.960 67.710 -10.860 ;
        RECT 65.410 -11.200 67.710 -10.960 ;
        RECT 65.410 -11.310 65.860 -11.200 ;
        RECT 67.260 -11.310 67.710 -11.200 ;
        RECT 68.920 -10.960 69.370 -10.860 ;
        RECT 69.760 -10.960 70.170 -10.530 ;
        RECT 72.920 -10.600 74.470 -10.380 ;
        RECT 74.850 -10.390 75.280 -10.330 ;
        RECT 75.660 -10.380 76.110 -10.330 ;
        RECT 76.710 -10.380 77.210 -9.990 ;
        RECT 75.660 -10.600 77.210 -10.380 ;
        RECT 86.420 -9.990 87.970 -9.770 ;
        RECT 86.420 -10.380 86.920 -9.990 ;
        RECT 87.520 -10.040 87.970 -9.990 ;
        RECT 88.350 -10.040 88.780 -9.980 ;
        RECT 89.160 -9.990 90.710 -9.770 ;
        RECT 93.460 -9.840 93.870 -9.410 ;
        RECT 94.260 -9.510 94.710 -9.410 ;
        RECT 95.920 -9.170 96.370 -9.060 ;
        RECT 97.770 -9.170 98.220 -9.060 ;
        RECT 95.920 -9.410 98.220 -9.170 ;
        RECT 95.920 -9.510 96.370 -9.410 ;
        RECT 96.760 -9.840 97.170 -9.410 ;
        RECT 97.770 -9.480 98.220 -9.410 ;
        RECT 99.170 -9.170 99.620 -9.090 ;
        RECT 100.220 -9.170 100.630 -8.730 ;
        RECT 101.020 -9.170 101.470 -9.060 ;
        RECT 99.170 -9.410 101.470 -9.170 ;
        RECT 99.170 -9.510 99.620 -9.410 ;
        RECT 101.020 -9.510 101.470 -9.410 ;
        RECT 102.660 -9.170 103.110 -9.060 ;
        RECT 103.500 -9.170 103.910 -8.730 ;
        RECT 106.680 -9.000 107.130 -8.720 ;
        RECT 110.500 -9.000 110.950 -8.720 ;
        RECT 120.180 -8.720 121.710 -8.510 ;
        RECT 122.090 -8.600 122.540 -8.510 ;
        RECT 122.920 -8.720 124.450 -8.510 ;
        RECT 104.510 -9.170 104.960 -9.090 ;
        RECT 102.660 -9.410 104.960 -9.170 ;
        RECT 102.660 -9.510 103.110 -9.410 ;
        RECT 104.510 -9.510 104.960 -9.410 ;
        RECT 105.910 -9.170 106.360 -9.060 ;
        RECT 107.760 -9.170 108.210 -9.060 ;
        RECT 105.910 -9.410 108.210 -9.170 ;
        RECT 105.910 -9.480 106.360 -9.410 ;
        RECT 89.160 -10.040 89.610 -9.990 ;
        RECT 87.520 -10.330 89.610 -10.040 ;
        RECT 87.520 -10.380 87.970 -10.330 ;
        RECT 70.770 -10.960 71.220 -10.890 ;
        RECT 68.920 -11.200 71.220 -10.960 ;
        RECT 68.920 -11.310 69.370 -11.200 ;
        RECT 70.770 -11.310 71.220 -11.200 ;
        RECT 72.170 -10.960 72.620 -10.860 ;
        RECT 74.020 -10.960 74.470 -10.860 ;
        RECT 72.170 -11.200 74.470 -10.960 ;
        RECT 72.170 -11.280 72.620 -11.200 ;
        RECT 52.680 -11.810 54.210 -11.650 ;
        RECT 54.590 -11.810 55.040 -11.770 ;
        RECT 55.420 -11.810 56.950 -11.650 ;
        RECT 52.680 -11.860 56.950 -11.810 ;
        RECT 66.180 -11.650 66.630 -11.370 ;
        RECT 70.000 -11.650 70.450 -11.370 ;
        RECT 73.220 -11.640 73.630 -11.200 ;
        RECT 74.020 -11.310 74.470 -11.200 ;
        RECT 75.660 -10.960 76.110 -10.860 ;
        RECT 77.510 -10.960 77.960 -10.860 ;
        RECT 75.660 -11.200 77.960 -10.960 ;
        RECT 75.660 -11.310 76.110 -11.200 ;
        RECT 76.500 -11.640 76.910 -11.200 ;
        RECT 77.510 -11.280 77.960 -11.200 ;
        RECT 78.910 -10.960 79.360 -10.890 ;
        RECT 79.960 -10.960 80.370 -10.530 ;
        RECT 80.760 -10.960 81.210 -10.860 ;
        RECT 78.910 -11.200 81.210 -10.960 ;
        RECT 78.910 -11.310 79.360 -11.200 ;
        RECT 80.760 -11.310 81.210 -11.200 ;
        RECT 82.420 -10.960 82.870 -10.860 ;
        RECT 83.260 -10.960 83.670 -10.530 ;
        RECT 86.420 -10.600 87.970 -10.380 ;
        RECT 88.350 -10.390 88.780 -10.330 ;
        RECT 89.160 -10.380 89.610 -10.330 ;
        RECT 90.210 -10.380 90.710 -9.990 ;
        RECT 89.160 -10.600 90.710 -10.380 ;
        RECT 99.920 -9.990 101.470 -9.770 ;
        RECT 99.920 -10.380 100.420 -9.990 ;
        RECT 101.020 -10.040 101.470 -9.990 ;
        RECT 101.850 -10.040 102.280 -9.980 ;
        RECT 102.660 -9.990 104.210 -9.770 ;
        RECT 106.960 -9.840 107.370 -9.410 ;
        RECT 107.760 -9.510 108.210 -9.410 ;
        RECT 109.420 -9.170 109.870 -9.060 ;
        RECT 111.270 -9.170 111.720 -9.060 ;
        RECT 109.420 -9.410 111.720 -9.170 ;
        RECT 109.420 -9.510 109.870 -9.410 ;
        RECT 110.260 -9.840 110.670 -9.410 ;
        RECT 111.270 -9.480 111.720 -9.410 ;
        RECT 112.670 -9.170 113.120 -9.090 ;
        RECT 113.720 -9.170 114.130 -8.730 ;
        RECT 114.520 -9.170 114.970 -9.060 ;
        RECT 112.670 -9.410 114.970 -9.170 ;
        RECT 112.670 -9.510 113.120 -9.410 ;
        RECT 114.520 -9.510 114.970 -9.410 ;
        RECT 116.160 -9.170 116.610 -9.060 ;
        RECT 117.000 -9.170 117.410 -8.730 ;
        RECT 120.180 -9.000 120.630 -8.720 ;
        RECT 124.000 -9.000 124.450 -8.720 ;
        RECT 133.680 -8.720 135.210 -8.510 ;
        RECT 135.590 -8.600 136.040 -8.510 ;
        RECT 136.420 -8.720 137.950 -8.510 ;
        RECT 118.010 -9.170 118.460 -9.090 ;
        RECT 116.160 -9.410 118.460 -9.170 ;
        RECT 116.160 -9.510 116.610 -9.410 ;
        RECT 118.010 -9.510 118.460 -9.410 ;
        RECT 119.410 -9.170 119.860 -9.060 ;
        RECT 121.260 -9.170 121.710 -9.060 ;
        RECT 119.410 -9.410 121.710 -9.170 ;
        RECT 119.410 -9.480 119.860 -9.410 ;
        RECT 102.660 -10.040 103.110 -9.990 ;
        RECT 101.020 -10.330 103.110 -10.040 ;
        RECT 101.020 -10.380 101.470 -10.330 ;
        RECT 84.270 -10.960 84.720 -10.890 ;
        RECT 82.420 -11.200 84.720 -10.960 ;
        RECT 82.420 -11.310 82.870 -11.200 ;
        RECT 84.270 -11.310 84.720 -11.200 ;
        RECT 85.670 -10.960 86.120 -10.860 ;
        RECT 87.520 -10.960 87.970 -10.860 ;
        RECT 85.670 -11.200 87.970 -10.960 ;
        RECT 85.670 -11.280 86.120 -11.200 ;
        RECT 66.180 -11.860 67.710 -11.650 ;
        RECT 68.090 -11.860 68.540 -11.770 ;
        RECT 68.920 -11.860 70.450 -11.650 ;
        RECT 79.680 -11.650 80.130 -11.370 ;
        RECT 83.500 -11.650 83.950 -11.370 ;
        RECT 86.720 -11.640 87.130 -11.200 ;
        RECT 87.520 -11.310 87.970 -11.200 ;
        RECT 89.160 -10.960 89.610 -10.860 ;
        RECT 91.010 -10.960 91.460 -10.860 ;
        RECT 89.160 -11.200 91.460 -10.960 ;
        RECT 89.160 -11.310 89.610 -11.200 ;
        RECT 90.000 -11.640 90.410 -11.200 ;
        RECT 91.010 -11.280 91.460 -11.200 ;
        RECT 92.410 -10.960 92.860 -10.890 ;
        RECT 93.460 -10.960 93.870 -10.530 ;
        RECT 94.260 -10.960 94.710 -10.860 ;
        RECT 92.410 -11.200 94.710 -10.960 ;
        RECT 92.410 -11.310 92.860 -11.200 ;
        RECT 94.260 -11.310 94.710 -11.200 ;
        RECT 95.920 -10.960 96.370 -10.860 ;
        RECT 96.760 -10.960 97.170 -10.530 ;
        RECT 99.920 -10.600 101.470 -10.380 ;
        RECT 101.850 -10.390 102.280 -10.330 ;
        RECT 102.660 -10.380 103.110 -10.330 ;
        RECT 103.710 -10.380 104.210 -9.990 ;
        RECT 102.660 -10.600 104.210 -10.380 ;
        RECT 113.420 -9.990 114.970 -9.770 ;
        RECT 113.420 -10.380 113.920 -9.990 ;
        RECT 114.520 -10.040 114.970 -9.990 ;
        RECT 115.350 -10.040 115.780 -9.980 ;
        RECT 116.160 -9.990 117.710 -9.770 ;
        RECT 120.460 -9.840 120.870 -9.410 ;
        RECT 121.260 -9.510 121.710 -9.410 ;
        RECT 122.920 -9.170 123.370 -9.060 ;
        RECT 124.770 -9.170 125.220 -9.060 ;
        RECT 122.920 -9.410 125.220 -9.170 ;
        RECT 122.920 -9.510 123.370 -9.410 ;
        RECT 123.760 -9.840 124.170 -9.410 ;
        RECT 124.770 -9.480 125.220 -9.410 ;
        RECT 126.170 -9.170 126.620 -9.090 ;
        RECT 127.220 -9.170 127.630 -8.730 ;
        RECT 128.020 -9.170 128.470 -9.060 ;
        RECT 126.170 -9.410 128.470 -9.170 ;
        RECT 126.170 -9.510 126.620 -9.410 ;
        RECT 128.020 -9.510 128.470 -9.410 ;
        RECT 129.660 -9.170 130.110 -9.060 ;
        RECT 130.500 -9.170 130.910 -8.730 ;
        RECT 133.680 -9.000 134.130 -8.720 ;
        RECT 137.500 -9.000 137.950 -8.720 ;
        RECT 147.180 -8.720 148.710 -8.510 ;
        RECT 149.090 -8.600 149.540 -8.510 ;
        RECT 149.920 -8.720 151.450 -8.510 ;
        RECT 131.510 -9.170 131.960 -9.090 ;
        RECT 129.660 -9.410 131.960 -9.170 ;
        RECT 129.660 -9.510 130.110 -9.410 ;
        RECT 131.510 -9.510 131.960 -9.410 ;
        RECT 132.910 -9.170 133.360 -9.060 ;
        RECT 134.760 -9.170 135.210 -9.060 ;
        RECT 132.910 -9.410 135.210 -9.170 ;
        RECT 132.910 -9.480 133.360 -9.410 ;
        RECT 116.160 -10.040 116.610 -9.990 ;
        RECT 114.520 -10.330 116.610 -10.040 ;
        RECT 114.520 -10.380 114.970 -10.330 ;
        RECT 97.770 -10.960 98.220 -10.890 ;
        RECT 95.920 -11.200 98.220 -10.960 ;
        RECT 95.920 -11.310 96.370 -11.200 ;
        RECT 97.770 -11.310 98.220 -11.200 ;
        RECT 99.170 -10.960 99.620 -10.860 ;
        RECT 101.020 -10.960 101.470 -10.860 ;
        RECT 99.170 -11.200 101.470 -10.960 ;
        RECT 99.170 -11.280 99.620 -11.200 ;
        RECT 79.680 -11.860 81.210 -11.650 ;
        RECT 81.590 -11.860 82.040 -11.770 ;
        RECT 82.420 -11.860 83.950 -11.650 ;
        RECT 93.180 -11.650 93.630 -11.370 ;
        RECT 97.000 -11.650 97.450 -11.370 ;
        RECT 100.220 -11.640 100.630 -11.200 ;
        RECT 101.020 -11.310 101.470 -11.200 ;
        RECT 102.660 -10.960 103.110 -10.860 ;
        RECT 104.510 -10.960 104.960 -10.860 ;
        RECT 102.660 -11.200 104.960 -10.960 ;
        RECT 102.660 -11.310 103.110 -11.200 ;
        RECT 103.500 -11.640 103.910 -11.200 ;
        RECT 104.510 -11.280 104.960 -11.200 ;
        RECT 105.910 -10.960 106.360 -10.890 ;
        RECT 106.960 -10.960 107.370 -10.530 ;
        RECT 107.760 -10.960 108.210 -10.860 ;
        RECT 105.910 -11.200 108.210 -10.960 ;
        RECT 105.910 -11.310 106.360 -11.200 ;
        RECT 107.760 -11.310 108.210 -11.200 ;
        RECT 109.420 -10.960 109.870 -10.860 ;
        RECT 110.260 -10.960 110.670 -10.530 ;
        RECT 113.420 -10.600 114.970 -10.380 ;
        RECT 115.350 -10.390 115.780 -10.330 ;
        RECT 116.160 -10.380 116.610 -10.330 ;
        RECT 117.210 -10.380 117.710 -9.990 ;
        RECT 116.160 -10.600 117.710 -10.380 ;
        RECT 126.920 -9.990 128.470 -9.770 ;
        RECT 126.920 -10.380 127.420 -9.990 ;
        RECT 128.020 -10.040 128.470 -9.990 ;
        RECT 128.850 -10.040 129.280 -9.980 ;
        RECT 129.660 -9.990 131.210 -9.770 ;
        RECT 133.960 -9.840 134.370 -9.410 ;
        RECT 134.760 -9.510 135.210 -9.410 ;
        RECT 136.420 -9.170 136.870 -9.060 ;
        RECT 138.270 -9.170 138.720 -9.060 ;
        RECT 136.420 -9.410 138.720 -9.170 ;
        RECT 136.420 -9.510 136.870 -9.410 ;
        RECT 137.260 -9.840 137.670 -9.410 ;
        RECT 138.270 -9.480 138.720 -9.410 ;
        RECT 139.670 -9.170 140.120 -9.090 ;
        RECT 140.720 -9.170 141.130 -8.730 ;
        RECT 141.520 -9.170 141.970 -9.060 ;
        RECT 139.670 -9.410 141.970 -9.170 ;
        RECT 139.670 -9.510 140.120 -9.410 ;
        RECT 141.520 -9.510 141.970 -9.410 ;
        RECT 143.160 -9.170 143.610 -9.060 ;
        RECT 144.000 -9.170 144.410 -8.730 ;
        RECT 147.180 -9.000 147.630 -8.720 ;
        RECT 151.000 -9.000 151.450 -8.720 ;
        RECT 160.680 -8.720 162.210 -8.510 ;
        RECT 162.590 -8.600 163.040 -8.510 ;
        RECT 163.420 -8.720 164.950 -8.510 ;
        RECT 145.010 -9.170 145.460 -9.090 ;
        RECT 143.160 -9.410 145.460 -9.170 ;
        RECT 143.160 -9.510 143.610 -9.410 ;
        RECT 145.010 -9.510 145.460 -9.410 ;
        RECT 146.410 -9.170 146.860 -9.060 ;
        RECT 148.260 -9.170 148.710 -9.060 ;
        RECT 146.410 -9.410 148.710 -9.170 ;
        RECT 146.410 -9.480 146.860 -9.410 ;
        RECT 129.660 -10.040 130.110 -9.990 ;
        RECT 128.020 -10.330 130.110 -10.040 ;
        RECT 128.020 -10.380 128.470 -10.330 ;
        RECT 111.270 -10.960 111.720 -10.890 ;
        RECT 109.420 -11.200 111.720 -10.960 ;
        RECT 109.420 -11.310 109.870 -11.200 ;
        RECT 111.270 -11.310 111.720 -11.200 ;
        RECT 112.670 -10.960 113.120 -10.860 ;
        RECT 114.520 -10.960 114.970 -10.860 ;
        RECT 112.670 -11.200 114.970 -10.960 ;
        RECT 112.670 -11.280 113.120 -11.200 ;
        RECT 93.180 -11.860 94.710 -11.650 ;
        RECT 95.090 -11.860 95.540 -11.770 ;
        RECT 95.920 -11.860 97.450 -11.650 ;
        RECT 106.680 -11.650 107.130 -11.370 ;
        RECT 110.500 -11.650 110.950 -11.370 ;
        RECT 113.720 -11.640 114.130 -11.200 ;
        RECT 114.520 -11.310 114.970 -11.200 ;
        RECT 116.160 -10.960 116.610 -10.860 ;
        RECT 118.010 -10.960 118.460 -10.860 ;
        RECT 116.160 -11.200 118.460 -10.960 ;
        RECT 116.160 -11.310 116.610 -11.200 ;
        RECT 117.000 -11.640 117.410 -11.200 ;
        RECT 118.010 -11.280 118.460 -11.200 ;
        RECT 119.410 -10.960 119.860 -10.890 ;
        RECT 120.460 -10.960 120.870 -10.530 ;
        RECT 121.260 -10.960 121.710 -10.860 ;
        RECT 119.410 -11.200 121.710 -10.960 ;
        RECT 119.410 -11.310 119.860 -11.200 ;
        RECT 121.260 -11.310 121.710 -11.200 ;
        RECT 122.920 -10.960 123.370 -10.860 ;
        RECT 123.760 -10.960 124.170 -10.530 ;
        RECT 126.920 -10.600 128.470 -10.380 ;
        RECT 128.850 -10.390 129.280 -10.330 ;
        RECT 129.660 -10.380 130.110 -10.330 ;
        RECT 130.710 -10.380 131.210 -9.990 ;
        RECT 129.660 -10.600 131.210 -10.380 ;
        RECT 140.420 -9.990 141.970 -9.770 ;
        RECT 140.420 -10.380 140.920 -9.990 ;
        RECT 141.520 -10.040 141.970 -9.990 ;
        RECT 142.350 -10.040 142.780 -9.980 ;
        RECT 143.160 -9.990 144.710 -9.770 ;
        RECT 147.460 -9.840 147.870 -9.410 ;
        RECT 148.260 -9.510 148.710 -9.410 ;
        RECT 149.920 -9.170 150.370 -9.060 ;
        RECT 151.770 -9.170 152.220 -9.060 ;
        RECT 149.920 -9.410 152.220 -9.170 ;
        RECT 149.920 -9.510 150.370 -9.410 ;
        RECT 150.760 -9.840 151.170 -9.410 ;
        RECT 151.770 -9.480 152.220 -9.410 ;
        RECT 153.170 -9.170 153.620 -9.090 ;
        RECT 154.220 -9.170 154.630 -8.730 ;
        RECT 155.020 -9.170 155.470 -9.060 ;
        RECT 153.170 -9.410 155.470 -9.170 ;
        RECT 153.170 -9.510 153.620 -9.410 ;
        RECT 155.020 -9.510 155.470 -9.410 ;
        RECT 156.660 -9.170 157.110 -9.060 ;
        RECT 157.500 -9.170 157.910 -8.730 ;
        RECT 160.680 -9.000 161.130 -8.720 ;
        RECT 164.500 -9.000 164.950 -8.720 ;
        RECT 174.180 -8.720 175.710 -8.510 ;
        RECT 176.090 -8.600 176.540 -8.510 ;
        RECT 176.920 -8.720 178.450 -8.510 ;
        RECT 158.510 -9.170 158.960 -9.090 ;
        RECT 156.660 -9.410 158.960 -9.170 ;
        RECT 156.660 -9.510 157.110 -9.410 ;
        RECT 158.510 -9.510 158.960 -9.410 ;
        RECT 159.910 -9.170 160.360 -9.060 ;
        RECT 161.760 -9.170 162.210 -9.060 ;
        RECT 159.910 -9.410 162.210 -9.170 ;
        RECT 159.910 -9.480 160.360 -9.410 ;
        RECT 143.160 -10.040 143.610 -9.990 ;
        RECT 141.520 -10.330 143.610 -10.040 ;
        RECT 141.520 -10.380 141.970 -10.330 ;
        RECT 124.770 -10.960 125.220 -10.890 ;
        RECT 122.920 -11.200 125.220 -10.960 ;
        RECT 122.920 -11.310 123.370 -11.200 ;
        RECT 124.770 -11.310 125.220 -11.200 ;
        RECT 126.170 -10.960 126.620 -10.860 ;
        RECT 128.020 -10.960 128.470 -10.860 ;
        RECT 126.170 -11.200 128.470 -10.960 ;
        RECT 126.170 -11.280 126.620 -11.200 ;
        RECT 106.680 -11.810 108.210 -11.650 ;
        RECT 108.590 -11.810 109.040 -11.770 ;
        RECT 109.420 -11.810 110.950 -11.650 ;
        RECT 106.680 -11.860 110.950 -11.810 ;
        RECT 120.180 -11.650 120.630 -11.370 ;
        RECT 124.000 -11.650 124.450 -11.370 ;
        RECT 127.220 -11.640 127.630 -11.200 ;
        RECT 128.020 -11.310 128.470 -11.200 ;
        RECT 129.660 -10.960 130.110 -10.860 ;
        RECT 131.510 -10.960 131.960 -10.860 ;
        RECT 129.660 -11.200 131.960 -10.960 ;
        RECT 129.660 -11.310 130.110 -11.200 ;
        RECT 130.500 -11.640 130.910 -11.200 ;
        RECT 131.510 -11.280 131.960 -11.200 ;
        RECT 132.910 -10.960 133.360 -10.890 ;
        RECT 133.960 -10.960 134.370 -10.530 ;
        RECT 134.760 -10.960 135.210 -10.860 ;
        RECT 132.910 -11.200 135.210 -10.960 ;
        RECT 132.910 -11.310 133.360 -11.200 ;
        RECT 134.760 -11.310 135.210 -11.200 ;
        RECT 136.420 -10.960 136.870 -10.860 ;
        RECT 137.260 -10.960 137.670 -10.530 ;
        RECT 140.420 -10.600 141.970 -10.380 ;
        RECT 142.350 -10.390 142.780 -10.330 ;
        RECT 143.160 -10.380 143.610 -10.330 ;
        RECT 144.210 -10.380 144.710 -9.990 ;
        RECT 143.160 -10.600 144.710 -10.380 ;
        RECT 153.920 -9.990 155.470 -9.770 ;
        RECT 153.920 -10.380 154.420 -9.990 ;
        RECT 155.020 -10.040 155.470 -9.990 ;
        RECT 155.850 -10.040 156.280 -9.980 ;
        RECT 156.660 -9.990 158.210 -9.770 ;
        RECT 160.960 -9.840 161.370 -9.410 ;
        RECT 161.760 -9.510 162.210 -9.410 ;
        RECT 163.420 -9.170 163.870 -9.060 ;
        RECT 165.270 -9.170 165.720 -9.060 ;
        RECT 163.420 -9.410 165.720 -9.170 ;
        RECT 163.420 -9.510 163.870 -9.410 ;
        RECT 164.260 -9.840 164.670 -9.410 ;
        RECT 165.270 -9.480 165.720 -9.410 ;
        RECT 166.670 -9.170 167.120 -9.090 ;
        RECT 167.720 -9.170 168.130 -8.730 ;
        RECT 168.520 -9.170 168.970 -9.060 ;
        RECT 166.670 -9.410 168.970 -9.170 ;
        RECT 166.670 -9.510 167.120 -9.410 ;
        RECT 168.520 -9.510 168.970 -9.410 ;
        RECT 170.160 -9.170 170.610 -9.060 ;
        RECT 171.000 -9.170 171.410 -8.730 ;
        RECT 174.180 -9.000 174.630 -8.720 ;
        RECT 178.000 -9.000 178.450 -8.720 ;
        RECT 187.680 -8.720 189.210 -8.510 ;
        RECT 189.590 -8.600 190.040 -8.510 ;
        RECT 190.420 -8.720 191.950 -8.510 ;
        RECT 172.010 -9.170 172.460 -9.090 ;
        RECT 170.160 -9.410 172.460 -9.170 ;
        RECT 170.160 -9.510 170.610 -9.410 ;
        RECT 172.010 -9.510 172.460 -9.410 ;
        RECT 173.410 -9.170 173.860 -9.060 ;
        RECT 175.260 -9.170 175.710 -9.060 ;
        RECT 173.410 -9.410 175.710 -9.170 ;
        RECT 173.410 -9.480 173.860 -9.410 ;
        RECT 156.660 -10.040 157.110 -9.990 ;
        RECT 155.020 -10.330 157.110 -10.040 ;
        RECT 155.020 -10.380 155.470 -10.330 ;
        RECT 138.270 -10.960 138.720 -10.890 ;
        RECT 136.420 -11.200 138.720 -10.960 ;
        RECT 136.420 -11.310 136.870 -11.200 ;
        RECT 138.270 -11.310 138.720 -11.200 ;
        RECT 139.670 -10.960 140.120 -10.860 ;
        RECT 141.520 -10.960 141.970 -10.860 ;
        RECT 139.670 -11.200 141.970 -10.960 ;
        RECT 139.670 -11.280 140.120 -11.200 ;
        RECT 120.180 -11.860 121.710 -11.650 ;
        RECT 122.090 -11.860 122.540 -11.770 ;
        RECT 122.920 -11.860 124.450 -11.650 ;
        RECT 133.680 -11.650 134.130 -11.370 ;
        RECT 137.500 -11.650 137.950 -11.370 ;
        RECT 140.720 -11.640 141.130 -11.200 ;
        RECT 141.520 -11.310 141.970 -11.200 ;
        RECT 143.160 -10.960 143.610 -10.860 ;
        RECT 145.010 -10.960 145.460 -10.860 ;
        RECT 143.160 -11.200 145.460 -10.960 ;
        RECT 143.160 -11.310 143.610 -11.200 ;
        RECT 144.000 -11.640 144.410 -11.200 ;
        RECT 145.010 -11.280 145.460 -11.200 ;
        RECT 146.410 -10.960 146.860 -10.890 ;
        RECT 147.460 -10.960 147.870 -10.530 ;
        RECT 148.260 -10.960 148.710 -10.860 ;
        RECT 146.410 -11.200 148.710 -10.960 ;
        RECT 146.410 -11.310 146.860 -11.200 ;
        RECT 148.260 -11.310 148.710 -11.200 ;
        RECT 149.920 -10.960 150.370 -10.860 ;
        RECT 150.760 -10.960 151.170 -10.530 ;
        RECT 153.920 -10.600 155.470 -10.380 ;
        RECT 155.850 -10.390 156.280 -10.330 ;
        RECT 156.660 -10.380 157.110 -10.330 ;
        RECT 157.710 -10.380 158.210 -9.990 ;
        RECT 156.660 -10.600 158.210 -10.380 ;
        RECT 167.420 -9.990 168.970 -9.770 ;
        RECT 167.420 -10.380 167.920 -9.990 ;
        RECT 168.520 -10.040 168.970 -9.990 ;
        RECT 169.350 -10.040 169.780 -9.980 ;
        RECT 170.160 -9.990 171.710 -9.770 ;
        RECT 174.460 -9.840 174.870 -9.410 ;
        RECT 175.260 -9.510 175.710 -9.410 ;
        RECT 176.920 -9.170 177.370 -9.060 ;
        RECT 178.770 -9.170 179.220 -9.060 ;
        RECT 176.920 -9.410 179.220 -9.170 ;
        RECT 176.920 -9.510 177.370 -9.410 ;
        RECT 177.760 -9.840 178.170 -9.410 ;
        RECT 178.770 -9.480 179.220 -9.410 ;
        RECT 180.170 -9.170 180.620 -9.090 ;
        RECT 181.220 -9.170 181.630 -8.730 ;
        RECT 182.020 -9.170 182.470 -9.060 ;
        RECT 180.170 -9.410 182.470 -9.170 ;
        RECT 180.170 -9.510 180.620 -9.410 ;
        RECT 182.020 -9.510 182.470 -9.410 ;
        RECT 183.660 -9.170 184.110 -9.060 ;
        RECT 184.500 -9.170 184.910 -8.730 ;
        RECT 187.680 -9.000 188.130 -8.720 ;
        RECT 191.500 -9.000 191.950 -8.720 ;
        RECT 201.180 -8.720 202.710 -8.510 ;
        RECT 203.090 -8.600 203.540 -8.510 ;
        RECT 203.920 -8.720 205.450 -8.510 ;
        RECT 185.510 -9.170 185.960 -9.090 ;
        RECT 183.660 -9.410 185.960 -9.170 ;
        RECT 183.660 -9.510 184.110 -9.410 ;
        RECT 185.510 -9.510 185.960 -9.410 ;
        RECT 186.910 -9.170 187.360 -9.060 ;
        RECT 188.760 -9.170 189.210 -9.060 ;
        RECT 186.910 -9.410 189.210 -9.170 ;
        RECT 186.910 -9.480 187.360 -9.410 ;
        RECT 170.160 -10.040 170.610 -9.990 ;
        RECT 168.520 -10.330 170.610 -10.040 ;
        RECT 168.520 -10.380 168.970 -10.330 ;
        RECT 151.770 -10.960 152.220 -10.890 ;
        RECT 149.920 -11.200 152.220 -10.960 ;
        RECT 149.920 -11.310 150.370 -11.200 ;
        RECT 151.770 -11.310 152.220 -11.200 ;
        RECT 153.170 -10.960 153.620 -10.860 ;
        RECT 155.020 -10.960 155.470 -10.860 ;
        RECT 153.170 -11.200 155.470 -10.960 ;
        RECT 153.170 -11.280 153.620 -11.200 ;
        RECT 133.680 -11.860 135.210 -11.650 ;
        RECT 135.590 -11.860 136.040 -11.770 ;
        RECT 136.420 -11.860 137.950 -11.650 ;
        RECT 147.180 -11.650 147.630 -11.370 ;
        RECT 151.000 -11.650 151.450 -11.370 ;
        RECT 154.220 -11.640 154.630 -11.200 ;
        RECT 155.020 -11.310 155.470 -11.200 ;
        RECT 156.660 -10.960 157.110 -10.860 ;
        RECT 158.510 -10.960 158.960 -10.860 ;
        RECT 156.660 -11.200 158.960 -10.960 ;
        RECT 156.660 -11.310 157.110 -11.200 ;
        RECT 157.500 -11.640 157.910 -11.200 ;
        RECT 158.510 -11.280 158.960 -11.200 ;
        RECT 159.910 -10.960 160.360 -10.890 ;
        RECT 160.960 -10.960 161.370 -10.530 ;
        RECT 161.760 -10.960 162.210 -10.860 ;
        RECT 159.910 -11.200 162.210 -10.960 ;
        RECT 159.910 -11.310 160.360 -11.200 ;
        RECT 161.760 -11.310 162.210 -11.200 ;
        RECT 163.420 -10.960 163.870 -10.860 ;
        RECT 164.260 -10.960 164.670 -10.530 ;
        RECT 167.420 -10.600 168.970 -10.380 ;
        RECT 169.350 -10.390 169.780 -10.330 ;
        RECT 170.160 -10.380 170.610 -10.330 ;
        RECT 171.210 -10.380 171.710 -9.990 ;
        RECT 170.160 -10.600 171.710 -10.380 ;
        RECT 180.920 -9.990 182.470 -9.770 ;
        RECT 180.920 -10.380 181.420 -9.990 ;
        RECT 182.020 -10.040 182.470 -9.990 ;
        RECT 182.850 -10.040 183.280 -9.980 ;
        RECT 183.660 -9.990 185.210 -9.770 ;
        RECT 187.960 -9.840 188.370 -9.410 ;
        RECT 188.760 -9.510 189.210 -9.410 ;
        RECT 190.420 -9.170 190.870 -9.060 ;
        RECT 192.270 -9.170 192.720 -9.060 ;
        RECT 190.420 -9.410 192.720 -9.170 ;
        RECT 190.420 -9.510 190.870 -9.410 ;
        RECT 191.260 -9.840 191.670 -9.410 ;
        RECT 192.270 -9.480 192.720 -9.410 ;
        RECT 193.670 -9.170 194.120 -9.090 ;
        RECT 194.720 -9.170 195.130 -8.730 ;
        RECT 195.520 -9.170 195.970 -9.060 ;
        RECT 193.670 -9.410 195.970 -9.170 ;
        RECT 193.670 -9.510 194.120 -9.410 ;
        RECT 195.520 -9.510 195.970 -9.410 ;
        RECT 197.160 -9.170 197.610 -9.060 ;
        RECT 198.000 -9.170 198.410 -8.730 ;
        RECT 201.180 -9.000 201.630 -8.720 ;
        RECT 205.000 -9.000 205.450 -8.720 ;
        RECT 214.680 -8.720 216.210 -8.510 ;
        RECT 216.590 -8.600 217.030 -8.510 ;
        RECT 199.010 -9.170 199.460 -9.090 ;
        RECT 197.160 -9.410 199.460 -9.170 ;
        RECT 197.160 -9.510 197.610 -9.410 ;
        RECT 199.010 -9.510 199.460 -9.410 ;
        RECT 200.410 -9.170 200.860 -9.060 ;
        RECT 202.260 -9.170 202.710 -9.060 ;
        RECT 200.410 -9.410 202.710 -9.170 ;
        RECT 200.410 -9.480 200.860 -9.410 ;
        RECT 183.660 -10.040 184.110 -9.990 ;
        RECT 182.020 -10.330 184.110 -10.040 ;
        RECT 182.020 -10.380 182.470 -10.330 ;
        RECT 165.270 -10.960 165.720 -10.890 ;
        RECT 163.420 -11.200 165.720 -10.960 ;
        RECT 163.420 -11.310 163.870 -11.200 ;
        RECT 165.270 -11.310 165.720 -11.200 ;
        RECT 166.670 -10.960 167.120 -10.860 ;
        RECT 168.520 -10.960 168.970 -10.860 ;
        RECT 166.670 -11.200 168.970 -10.960 ;
        RECT 166.670 -11.280 167.120 -11.200 ;
        RECT 147.180 -11.860 148.710 -11.650 ;
        RECT 149.090 -11.860 149.540 -11.770 ;
        RECT 149.920 -11.860 151.450 -11.650 ;
        RECT 160.680 -11.650 161.130 -11.370 ;
        RECT 164.500 -11.650 164.950 -11.370 ;
        RECT 167.720 -11.640 168.130 -11.200 ;
        RECT 168.520 -11.310 168.970 -11.200 ;
        RECT 170.160 -10.960 170.610 -10.860 ;
        RECT 172.010 -10.960 172.460 -10.860 ;
        RECT 170.160 -11.200 172.460 -10.960 ;
        RECT 170.160 -11.310 170.610 -11.200 ;
        RECT 171.000 -11.640 171.410 -11.200 ;
        RECT 172.010 -11.280 172.460 -11.200 ;
        RECT 173.410 -10.960 173.860 -10.890 ;
        RECT 174.460 -10.960 174.870 -10.530 ;
        RECT 175.260 -10.960 175.710 -10.860 ;
        RECT 173.410 -11.200 175.710 -10.960 ;
        RECT 173.410 -11.310 173.860 -11.200 ;
        RECT 175.260 -11.310 175.710 -11.200 ;
        RECT 176.920 -10.960 177.370 -10.860 ;
        RECT 177.760 -10.960 178.170 -10.530 ;
        RECT 180.920 -10.600 182.470 -10.380 ;
        RECT 182.850 -10.390 183.280 -10.330 ;
        RECT 183.660 -10.380 184.110 -10.330 ;
        RECT 184.710 -10.380 185.210 -9.990 ;
        RECT 183.660 -10.600 185.210 -10.380 ;
        RECT 194.420 -9.990 195.970 -9.770 ;
        RECT 194.420 -10.380 194.920 -9.990 ;
        RECT 195.520 -10.040 195.970 -9.990 ;
        RECT 196.350 -10.040 196.780 -9.980 ;
        RECT 197.160 -9.990 198.710 -9.770 ;
        RECT 201.460 -9.840 201.870 -9.410 ;
        RECT 202.260 -9.510 202.710 -9.410 ;
        RECT 203.920 -9.170 204.370 -9.060 ;
        RECT 205.770 -9.170 206.220 -9.060 ;
        RECT 203.920 -9.410 206.220 -9.170 ;
        RECT 203.920 -9.510 204.370 -9.410 ;
        RECT 204.760 -9.840 205.170 -9.410 ;
        RECT 205.770 -9.480 206.220 -9.410 ;
        RECT 207.170 -9.170 207.620 -9.090 ;
        RECT 208.220 -9.170 208.630 -8.730 ;
        RECT 209.020 -9.170 209.470 -9.060 ;
        RECT 207.170 -9.410 209.470 -9.170 ;
        RECT 207.170 -9.510 207.620 -9.410 ;
        RECT 209.020 -9.510 209.470 -9.410 ;
        RECT 210.660 -9.170 211.110 -9.060 ;
        RECT 211.500 -9.170 211.910 -8.730 ;
        RECT 214.680 -9.000 215.130 -8.720 ;
        RECT 212.510 -9.170 212.960 -9.090 ;
        RECT 210.660 -9.410 212.960 -9.170 ;
        RECT 210.660 -9.510 211.110 -9.410 ;
        RECT 212.510 -9.510 212.960 -9.410 ;
        RECT 213.910 -9.170 214.360 -9.060 ;
        RECT 215.760 -9.170 216.210 -9.060 ;
        RECT 213.910 -9.410 216.210 -9.170 ;
        RECT 213.910 -9.480 214.360 -9.410 ;
        RECT 197.160 -10.040 197.610 -9.990 ;
        RECT 195.520 -10.330 197.610 -10.040 ;
        RECT 195.520 -10.380 195.970 -10.330 ;
        RECT 178.770 -10.960 179.220 -10.890 ;
        RECT 176.920 -11.200 179.220 -10.960 ;
        RECT 176.920 -11.310 177.370 -11.200 ;
        RECT 178.770 -11.310 179.220 -11.200 ;
        RECT 180.170 -10.960 180.620 -10.860 ;
        RECT 182.020 -10.960 182.470 -10.860 ;
        RECT 180.170 -11.200 182.470 -10.960 ;
        RECT 180.170 -11.280 180.620 -11.200 ;
        RECT 160.680 -11.810 162.210 -11.650 ;
        RECT 162.590 -11.810 163.040 -11.770 ;
        RECT 163.420 -11.810 164.950 -11.650 ;
        RECT 160.680 -11.860 164.950 -11.810 ;
        RECT 174.180 -11.650 174.630 -11.370 ;
        RECT 178.000 -11.650 178.450 -11.370 ;
        RECT 181.220 -11.640 181.630 -11.200 ;
        RECT 182.020 -11.310 182.470 -11.200 ;
        RECT 183.660 -10.960 184.110 -10.860 ;
        RECT 185.510 -10.960 185.960 -10.860 ;
        RECT 183.660 -11.200 185.960 -10.960 ;
        RECT 183.660 -11.310 184.110 -11.200 ;
        RECT 184.500 -11.640 184.910 -11.200 ;
        RECT 185.510 -11.280 185.960 -11.200 ;
        RECT 186.910 -10.960 187.360 -10.890 ;
        RECT 187.960 -10.960 188.370 -10.530 ;
        RECT 188.760 -10.960 189.210 -10.860 ;
        RECT 186.910 -11.200 189.210 -10.960 ;
        RECT 186.910 -11.310 187.360 -11.200 ;
        RECT 188.760 -11.310 189.210 -11.200 ;
        RECT 190.420 -10.960 190.870 -10.860 ;
        RECT 191.260 -10.960 191.670 -10.530 ;
        RECT 194.420 -10.600 195.970 -10.380 ;
        RECT 196.350 -10.390 196.780 -10.330 ;
        RECT 197.160 -10.380 197.610 -10.330 ;
        RECT 198.210 -10.380 198.710 -9.990 ;
        RECT 197.160 -10.600 198.710 -10.380 ;
        RECT 207.920 -9.990 209.470 -9.770 ;
        RECT 207.920 -10.380 208.420 -9.990 ;
        RECT 209.020 -10.040 209.470 -9.990 ;
        RECT 209.850 -10.040 210.280 -9.980 ;
        RECT 210.660 -9.990 212.210 -9.770 ;
        RECT 214.960 -9.840 215.370 -9.410 ;
        RECT 215.760 -9.510 216.210 -9.410 ;
        RECT 210.660 -10.040 211.110 -9.990 ;
        RECT 209.020 -10.330 211.110 -10.040 ;
        RECT 209.020 -10.380 209.470 -10.330 ;
        RECT 192.270 -10.960 192.720 -10.890 ;
        RECT 190.420 -11.200 192.720 -10.960 ;
        RECT 190.420 -11.310 190.870 -11.200 ;
        RECT 192.270 -11.310 192.720 -11.200 ;
        RECT 193.670 -10.960 194.120 -10.860 ;
        RECT 195.520 -10.960 195.970 -10.860 ;
        RECT 193.670 -11.200 195.970 -10.960 ;
        RECT 193.670 -11.280 194.120 -11.200 ;
        RECT 174.180 -11.860 175.710 -11.650 ;
        RECT 176.090 -11.860 176.540 -11.770 ;
        RECT 176.920 -11.860 178.450 -11.650 ;
        RECT 187.680 -11.650 188.130 -11.370 ;
        RECT 191.500 -11.650 191.950 -11.370 ;
        RECT 194.720 -11.640 195.130 -11.200 ;
        RECT 195.520 -11.310 195.970 -11.200 ;
        RECT 197.160 -10.960 197.610 -10.860 ;
        RECT 199.010 -10.960 199.460 -10.860 ;
        RECT 197.160 -11.200 199.460 -10.960 ;
        RECT 197.160 -11.310 197.610 -11.200 ;
        RECT 198.000 -11.640 198.410 -11.200 ;
        RECT 199.010 -11.280 199.460 -11.200 ;
        RECT 200.410 -10.960 200.860 -10.890 ;
        RECT 201.460 -10.960 201.870 -10.530 ;
        RECT 202.260 -10.960 202.710 -10.860 ;
        RECT 200.410 -11.200 202.710 -10.960 ;
        RECT 200.410 -11.310 200.860 -11.200 ;
        RECT 202.260 -11.310 202.710 -11.200 ;
        RECT 203.920 -10.960 204.370 -10.860 ;
        RECT 204.760 -10.960 205.170 -10.530 ;
        RECT 207.920 -10.600 209.470 -10.380 ;
        RECT 209.850 -10.390 210.280 -10.330 ;
        RECT 210.660 -10.380 211.110 -10.330 ;
        RECT 211.710 -10.380 212.210 -9.990 ;
        RECT 210.660 -10.600 212.210 -10.380 ;
        RECT 205.770 -10.960 206.220 -10.890 ;
        RECT 203.920 -11.200 206.220 -10.960 ;
        RECT 203.920 -11.310 204.370 -11.200 ;
        RECT 205.770 -11.310 206.220 -11.200 ;
        RECT 207.170 -10.960 207.620 -10.860 ;
        RECT 209.020 -10.960 209.470 -10.860 ;
        RECT 207.170 -11.200 209.470 -10.960 ;
        RECT 207.170 -11.280 207.620 -11.200 ;
        RECT 187.680 -11.860 189.210 -11.650 ;
        RECT 189.590 -11.860 190.040 -11.770 ;
        RECT 190.420 -11.860 191.950 -11.650 ;
        RECT 201.180 -11.650 201.630 -11.370 ;
        RECT 205.000 -11.650 205.450 -11.370 ;
        RECT 208.220 -11.640 208.630 -11.200 ;
        RECT 209.020 -11.310 209.470 -11.200 ;
        RECT 210.660 -10.960 211.110 -10.860 ;
        RECT 212.510 -10.960 212.960 -10.860 ;
        RECT 210.660 -11.200 212.960 -10.960 ;
        RECT 210.660 -11.310 211.110 -11.200 ;
        RECT 211.500 -11.640 211.910 -11.200 ;
        RECT 212.510 -11.280 212.960 -11.200 ;
        RECT 213.910 -10.960 214.360 -10.890 ;
        RECT 214.960 -10.960 215.370 -10.530 ;
        RECT 215.760 -10.960 216.210 -10.860 ;
        RECT 213.910 -11.200 216.210 -10.960 ;
        RECT 213.910 -11.310 214.360 -11.200 ;
        RECT 215.760 -11.310 216.210 -11.200 ;
        RECT 201.180 -11.860 202.710 -11.650 ;
        RECT 203.090 -11.860 203.540 -11.770 ;
        RECT 203.920 -11.860 205.450 -11.650 ;
        RECT 214.680 -11.650 215.130 -11.370 ;
        RECT 214.680 -11.860 216.210 -11.650 ;
        RECT 216.590 -11.810 217.030 -11.770 ;
        RECT 216.590 -11.860 217.690 -11.810 ;
        RECT 13.260 -12.120 15.370 -11.860 ;
        RECT 26.760 -12.120 28.870 -11.860 ;
        RECT 40.260 -12.120 42.370 -11.860 ;
        RECT 53.760 -12.120 55.870 -11.860 ;
        RECT 67.260 -12.120 69.370 -11.860 ;
        RECT 80.760 -12.120 82.870 -11.860 ;
        RECT 94.260 -12.120 96.370 -11.860 ;
        RECT 107.760 -12.120 109.870 -11.860 ;
        RECT 121.260 -12.120 123.370 -11.860 ;
        RECT 134.760 -12.120 136.870 -11.860 ;
        RECT 148.260 -12.120 150.370 -11.860 ;
        RECT 161.760 -12.120 163.870 -11.860 ;
        RECT 175.260 -12.120 177.370 -11.860 ;
        RECT 188.760 -12.120 190.870 -11.860 ;
        RECT 202.260 -12.120 204.370 -11.860 ;
        RECT 215.760 -12.120 217.690 -11.860 ;
        RECT 12.180 -12.330 13.710 -12.120 ;
        RECT 14.090 -12.210 14.540 -12.120 ;
        RECT 14.920 -12.330 16.450 -12.120 ;
        RECT 1.420 -12.780 1.870 -12.670 ;
        RECT 3.270 -12.780 3.720 -12.670 ;
        RECT 1.420 -13.020 3.720 -12.780 ;
        RECT 1.420 -13.120 1.870 -13.020 ;
        RECT 2.260 -13.450 2.670 -13.020 ;
        RECT 3.270 -13.090 3.720 -13.020 ;
        RECT 4.670 -12.780 5.120 -12.700 ;
        RECT 5.720 -12.780 6.130 -12.340 ;
        RECT 6.520 -12.780 6.970 -12.670 ;
        RECT 4.670 -13.020 6.970 -12.780 ;
        RECT 4.670 -13.120 5.120 -13.020 ;
        RECT 6.520 -13.120 6.970 -13.020 ;
        RECT 8.160 -12.780 8.610 -12.670 ;
        RECT 9.000 -12.780 9.410 -12.340 ;
        RECT 12.180 -12.610 12.630 -12.330 ;
        RECT 16.000 -12.610 16.450 -12.330 ;
        RECT 25.680 -12.330 27.210 -12.120 ;
        RECT 27.590 -12.210 28.040 -12.120 ;
        RECT 28.420 -12.330 29.950 -12.120 ;
        RECT 10.010 -12.780 10.460 -12.700 ;
        RECT 8.160 -13.020 10.460 -12.780 ;
        RECT 8.160 -13.120 8.610 -13.020 ;
        RECT 10.010 -13.120 10.460 -13.020 ;
        RECT 11.410 -12.780 11.860 -12.670 ;
        RECT 13.260 -12.780 13.710 -12.670 ;
        RECT 11.410 -13.020 13.710 -12.780 ;
        RECT 11.410 -13.090 11.860 -13.020 ;
        RECT 5.420 -13.600 6.970 -13.380 ;
        RECT 5.420 -13.990 5.920 -13.600 ;
        RECT 6.520 -13.650 6.970 -13.600 ;
        RECT 7.350 -13.650 7.780 -13.590 ;
        RECT 8.160 -13.600 9.710 -13.380 ;
        RECT 12.460 -13.450 12.870 -13.020 ;
        RECT 13.260 -13.120 13.710 -13.020 ;
        RECT 14.920 -12.780 15.370 -12.670 ;
        RECT 16.770 -12.780 17.220 -12.670 ;
        RECT 14.920 -13.020 17.220 -12.780 ;
        RECT 14.920 -13.120 15.370 -13.020 ;
        RECT 15.760 -13.450 16.170 -13.020 ;
        RECT 16.770 -13.090 17.220 -13.020 ;
        RECT 18.170 -12.780 18.620 -12.700 ;
        RECT 19.220 -12.780 19.630 -12.340 ;
        RECT 20.020 -12.780 20.470 -12.670 ;
        RECT 18.170 -13.020 20.470 -12.780 ;
        RECT 18.170 -13.120 18.620 -13.020 ;
        RECT 20.020 -13.120 20.470 -13.020 ;
        RECT 21.660 -12.780 22.110 -12.670 ;
        RECT 22.500 -12.780 22.910 -12.340 ;
        RECT 25.680 -12.610 26.130 -12.330 ;
        RECT 29.500 -12.610 29.950 -12.330 ;
        RECT 39.180 -12.330 40.710 -12.120 ;
        RECT 41.090 -12.210 41.540 -12.120 ;
        RECT 41.920 -12.330 43.450 -12.120 ;
        RECT 23.510 -12.780 23.960 -12.700 ;
        RECT 21.660 -13.020 23.960 -12.780 ;
        RECT 21.660 -13.120 22.110 -13.020 ;
        RECT 23.510 -13.120 23.960 -13.020 ;
        RECT 24.910 -12.780 25.360 -12.670 ;
        RECT 26.760 -12.780 27.210 -12.670 ;
        RECT 24.910 -13.020 27.210 -12.780 ;
        RECT 24.910 -13.090 25.360 -13.020 ;
        RECT 8.160 -13.650 8.610 -13.600 ;
        RECT 6.520 -13.940 8.610 -13.650 ;
        RECT 6.520 -13.990 6.970 -13.940 ;
        RECT 1.420 -14.570 1.870 -14.470 ;
        RECT 2.260 -14.570 2.670 -14.140 ;
        RECT 5.420 -14.210 6.970 -13.990 ;
        RECT 7.350 -14.000 7.780 -13.940 ;
        RECT 8.160 -13.990 8.610 -13.940 ;
        RECT 9.210 -13.990 9.710 -13.600 ;
        RECT 8.160 -14.210 9.710 -13.990 ;
        RECT 18.920 -13.600 20.470 -13.380 ;
        RECT 18.920 -13.990 19.420 -13.600 ;
        RECT 20.020 -13.650 20.470 -13.600 ;
        RECT 20.850 -13.650 21.280 -13.590 ;
        RECT 21.660 -13.600 23.210 -13.380 ;
        RECT 25.960 -13.450 26.370 -13.020 ;
        RECT 26.760 -13.120 27.210 -13.020 ;
        RECT 28.420 -12.780 28.870 -12.670 ;
        RECT 30.270 -12.780 30.720 -12.670 ;
        RECT 28.420 -13.020 30.720 -12.780 ;
        RECT 28.420 -13.120 28.870 -13.020 ;
        RECT 29.260 -13.450 29.670 -13.020 ;
        RECT 30.270 -13.090 30.720 -13.020 ;
        RECT 31.670 -12.780 32.120 -12.700 ;
        RECT 32.720 -12.780 33.130 -12.340 ;
        RECT 33.520 -12.780 33.970 -12.670 ;
        RECT 31.670 -13.020 33.970 -12.780 ;
        RECT 31.670 -13.120 32.120 -13.020 ;
        RECT 33.520 -13.120 33.970 -13.020 ;
        RECT 35.160 -12.780 35.610 -12.670 ;
        RECT 36.000 -12.780 36.410 -12.340 ;
        RECT 39.180 -12.610 39.630 -12.330 ;
        RECT 43.000 -12.610 43.450 -12.330 ;
        RECT 52.680 -12.170 56.950 -12.120 ;
        RECT 52.680 -12.330 54.210 -12.170 ;
        RECT 54.590 -12.210 55.040 -12.170 ;
        RECT 55.420 -12.330 56.950 -12.170 ;
        RECT 37.010 -12.780 37.460 -12.700 ;
        RECT 35.160 -13.020 37.460 -12.780 ;
        RECT 35.160 -13.120 35.610 -13.020 ;
        RECT 37.010 -13.120 37.460 -13.020 ;
        RECT 38.410 -12.780 38.860 -12.670 ;
        RECT 40.260 -12.780 40.710 -12.670 ;
        RECT 38.410 -13.020 40.710 -12.780 ;
        RECT 38.410 -13.090 38.860 -13.020 ;
        RECT 21.660 -13.650 22.110 -13.600 ;
        RECT 20.020 -13.940 22.110 -13.650 ;
        RECT 20.020 -13.990 20.470 -13.940 ;
        RECT 3.270 -14.570 3.720 -14.500 ;
        RECT 1.420 -14.810 3.720 -14.570 ;
        RECT 1.420 -14.920 1.870 -14.810 ;
        RECT 3.270 -14.920 3.720 -14.810 ;
        RECT 4.670 -14.570 5.120 -14.470 ;
        RECT 6.520 -14.570 6.970 -14.470 ;
        RECT 4.670 -14.810 6.970 -14.570 ;
        RECT 4.670 -14.890 5.120 -14.810 ;
        RECT 5.720 -15.250 6.130 -14.810 ;
        RECT 6.520 -14.920 6.970 -14.810 ;
        RECT 8.160 -14.570 8.610 -14.470 ;
        RECT 10.010 -14.570 10.460 -14.470 ;
        RECT 8.160 -14.810 10.460 -14.570 ;
        RECT 8.160 -14.920 8.610 -14.810 ;
        RECT 9.000 -15.250 9.410 -14.810 ;
        RECT 10.010 -14.890 10.460 -14.810 ;
        RECT 11.410 -14.570 11.860 -14.500 ;
        RECT 12.460 -14.570 12.870 -14.140 ;
        RECT 13.260 -14.570 13.710 -14.470 ;
        RECT 11.410 -14.810 13.710 -14.570 ;
        RECT 11.410 -14.920 11.860 -14.810 ;
        RECT 13.260 -14.920 13.710 -14.810 ;
        RECT 14.920 -14.570 15.370 -14.470 ;
        RECT 15.760 -14.570 16.170 -14.140 ;
        RECT 18.920 -14.210 20.470 -13.990 ;
        RECT 20.850 -14.000 21.280 -13.940 ;
        RECT 21.660 -13.990 22.110 -13.940 ;
        RECT 22.710 -13.990 23.210 -13.600 ;
        RECT 21.660 -14.210 23.210 -13.990 ;
        RECT 32.420 -13.600 33.970 -13.380 ;
        RECT 32.420 -13.990 32.920 -13.600 ;
        RECT 33.520 -13.650 33.970 -13.600 ;
        RECT 34.350 -13.650 34.780 -13.590 ;
        RECT 35.160 -13.600 36.710 -13.380 ;
        RECT 39.460 -13.450 39.870 -13.020 ;
        RECT 40.260 -13.120 40.710 -13.020 ;
        RECT 41.920 -12.780 42.370 -12.670 ;
        RECT 43.770 -12.780 44.220 -12.670 ;
        RECT 41.920 -13.020 44.220 -12.780 ;
        RECT 41.920 -13.120 42.370 -13.020 ;
        RECT 42.760 -13.450 43.170 -13.020 ;
        RECT 43.770 -13.090 44.220 -13.020 ;
        RECT 45.170 -12.780 45.620 -12.700 ;
        RECT 46.220 -12.780 46.630 -12.340 ;
        RECT 47.020 -12.780 47.470 -12.670 ;
        RECT 45.170 -13.020 47.470 -12.780 ;
        RECT 45.170 -13.120 45.620 -13.020 ;
        RECT 47.020 -13.120 47.470 -13.020 ;
        RECT 48.660 -12.780 49.110 -12.670 ;
        RECT 49.500 -12.780 49.910 -12.340 ;
        RECT 52.680 -12.610 53.130 -12.330 ;
        RECT 56.500 -12.610 56.950 -12.330 ;
        RECT 66.180 -12.330 67.710 -12.120 ;
        RECT 68.090 -12.210 68.540 -12.120 ;
        RECT 68.920 -12.330 70.450 -12.120 ;
        RECT 50.510 -12.780 50.960 -12.700 ;
        RECT 48.660 -13.020 50.960 -12.780 ;
        RECT 48.660 -13.120 49.110 -13.020 ;
        RECT 50.510 -13.120 50.960 -13.020 ;
        RECT 51.910 -12.780 52.360 -12.670 ;
        RECT 53.760 -12.780 54.210 -12.670 ;
        RECT 51.910 -13.020 54.210 -12.780 ;
        RECT 51.910 -13.090 52.360 -13.020 ;
        RECT 35.160 -13.650 35.610 -13.600 ;
        RECT 33.520 -13.940 35.610 -13.650 ;
        RECT 33.520 -13.990 33.970 -13.940 ;
        RECT 16.770 -14.570 17.220 -14.500 ;
        RECT 14.920 -14.810 17.220 -14.570 ;
        RECT 14.920 -14.920 15.370 -14.810 ;
        RECT 16.770 -14.920 17.220 -14.810 ;
        RECT 18.170 -14.570 18.620 -14.470 ;
        RECT 20.020 -14.570 20.470 -14.470 ;
        RECT 18.170 -14.810 20.470 -14.570 ;
        RECT 18.170 -14.890 18.620 -14.810 ;
        RECT 12.180 -15.260 12.630 -14.980 ;
        RECT 16.000 -15.260 16.450 -14.980 ;
        RECT 19.220 -15.250 19.630 -14.810 ;
        RECT 20.020 -14.920 20.470 -14.810 ;
        RECT 21.660 -14.570 22.110 -14.470 ;
        RECT 23.510 -14.570 23.960 -14.470 ;
        RECT 21.660 -14.810 23.960 -14.570 ;
        RECT 21.660 -14.920 22.110 -14.810 ;
        RECT 22.500 -15.250 22.910 -14.810 ;
        RECT 23.510 -14.890 23.960 -14.810 ;
        RECT 24.910 -14.570 25.360 -14.500 ;
        RECT 25.960 -14.570 26.370 -14.140 ;
        RECT 26.760 -14.570 27.210 -14.470 ;
        RECT 24.910 -14.810 27.210 -14.570 ;
        RECT 24.910 -14.920 25.360 -14.810 ;
        RECT 26.760 -14.920 27.210 -14.810 ;
        RECT 28.420 -14.570 28.870 -14.470 ;
        RECT 29.260 -14.570 29.670 -14.140 ;
        RECT 32.420 -14.210 33.970 -13.990 ;
        RECT 34.350 -14.000 34.780 -13.940 ;
        RECT 35.160 -13.990 35.610 -13.940 ;
        RECT 36.210 -13.990 36.710 -13.600 ;
        RECT 35.160 -14.210 36.710 -13.990 ;
        RECT 45.920 -13.600 47.470 -13.380 ;
        RECT 45.920 -13.990 46.420 -13.600 ;
        RECT 47.020 -13.650 47.470 -13.600 ;
        RECT 47.850 -13.650 48.280 -13.590 ;
        RECT 48.660 -13.600 50.210 -13.380 ;
        RECT 52.960 -13.450 53.370 -13.020 ;
        RECT 53.760 -13.120 54.210 -13.020 ;
        RECT 55.420 -12.780 55.870 -12.670 ;
        RECT 57.270 -12.780 57.720 -12.670 ;
        RECT 55.420 -13.020 57.720 -12.780 ;
        RECT 55.420 -13.120 55.870 -13.020 ;
        RECT 56.260 -13.450 56.670 -13.020 ;
        RECT 57.270 -13.090 57.720 -13.020 ;
        RECT 58.670 -12.780 59.120 -12.700 ;
        RECT 59.720 -12.780 60.130 -12.340 ;
        RECT 60.520 -12.780 60.970 -12.670 ;
        RECT 58.670 -13.020 60.970 -12.780 ;
        RECT 58.670 -13.120 59.120 -13.020 ;
        RECT 60.520 -13.120 60.970 -13.020 ;
        RECT 62.160 -12.780 62.610 -12.670 ;
        RECT 63.000 -12.780 63.410 -12.340 ;
        RECT 66.180 -12.610 66.630 -12.330 ;
        RECT 70.000 -12.610 70.450 -12.330 ;
        RECT 79.680 -12.330 81.210 -12.120 ;
        RECT 81.590 -12.210 82.040 -12.120 ;
        RECT 82.420 -12.330 83.950 -12.120 ;
        RECT 64.010 -12.780 64.460 -12.700 ;
        RECT 62.160 -13.020 64.460 -12.780 ;
        RECT 62.160 -13.120 62.610 -13.020 ;
        RECT 64.010 -13.120 64.460 -13.020 ;
        RECT 65.410 -12.780 65.860 -12.670 ;
        RECT 67.260 -12.780 67.710 -12.670 ;
        RECT 65.410 -13.020 67.710 -12.780 ;
        RECT 65.410 -13.090 65.860 -13.020 ;
        RECT 48.660 -13.650 49.110 -13.600 ;
        RECT 47.020 -13.940 49.110 -13.650 ;
        RECT 47.020 -13.990 47.470 -13.940 ;
        RECT 30.270 -14.570 30.720 -14.500 ;
        RECT 28.420 -14.810 30.720 -14.570 ;
        RECT 28.420 -14.920 28.870 -14.810 ;
        RECT 30.270 -14.920 30.720 -14.810 ;
        RECT 31.670 -14.570 32.120 -14.470 ;
        RECT 33.520 -14.570 33.970 -14.470 ;
        RECT 31.670 -14.810 33.970 -14.570 ;
        RECT 31.670 -14.890 32.120 -14.810 ;
        RECT 12.180 -15.470 13.710 -15.260 ;
        RECT 14.090 -15.470 14.540 -15.380 ;
        RECT 14.920 -15.470 16.450 -15.260 ;
        RECT 25.680 -15.260 26.130 -14.980 ;
        RECT 29.500 -15.260 29.950 -14.980 ;
        RECT 32.720 -15.250 33.130 -14.810 ;
        RECT 33.520 -14.920 33.970 -14.810 ;
        RECT 35.160 -14.570 35.610 -14.470 ;
        RECT 37.010 -14.570 37.460 -14.470 ;
        RECT 35.160 -14.810 37.460 -14.570 ;
        RECT 35.160 -14.920 35.610 -14.810 ;
        RECT 36.000 -15.250 36.410 -14.810 ;
        RECT 37.010 -14.890 37.460 -14.810 ;
        RECT 38.410 -14.570 38.860 -14.500 ;
        RECT 39.460 -14.570 39.870 -14.140 ;
        RECT 40.260 -14.570 40.710 -14.470 ;
        RECT 38.410 -14.810 40.710 -14.570 ;
        RECT 38.410 -14.920 38.860 -14.810 ;
        RECT 40.260 -14.920 40.710 -14.810 ;
        RECT 41.920 -14.570 42.370 -14.470 ;
        RECT 42.760 -14.570 43.170 -14.140 ;
        RECT 45.920 -14.210 47.470 -13.990 ;
        RECT 47.850 -14.000 48.280 -13.940 ;
        RECT 48.660 -13.990 49.110 -13.940 ;
        RECT 49.710 -13.990 50.210 -13.600 ;
        RECT 48.660 -14.210 50.210 -13.990 ;
        RECT 59.420 -13.600 60.970 -13.380 ;
        RECT 59.420 -13.990 59.920 -13.600 ;
        RECT 60.520 -13.650 60.970 -13.600 ;
        RECT 61.350 -13.650 61.780 -13.590 ;
        RECT 62.160 -13.600 63.710 -13.380 ;
        RECT 66.460 -13.450 66.870 -13.020 ;
        RECT 67.260 -13.120 67.710 -13.020 ;
        RECT 68.920 -12.780 69.370 -12.670 ;
        RECT 70.770 -12.780 71.220 -12.670 ;
        RECT 68.920 -13.020 71.220 -12.780 ;
        RECT 68.920 -13.120 69.370 -13.020 ;
        RECT 69.760 -13.450 70.170 -13.020 ;
        RECT 70.770 -13.090 71.220 -13.020 ;
        RECT 72.170 -12.780 72.620 -12.700 ;
        RECT 73.220 -12.780 73.630 -12.340 ;
        RECT 74.020 -12.780 74.470 -12.670 ;
        RECT 72.170 -13.020 74.470 -12.780 ;
        RECT 72.170 -13.120 72.620 -13.020 ;
        RECT 74.020 -13.120 74.470 -13.020 ;
        RECT 75.660 -12.780 76.110 -12.670 ;
        RECT 76.500 -12.780 76.910 -12.340 ;
        RECT 79.680 -12.610 80.130 -12.330 ;
        RECT 83.500 -12.610 83.950 -12.330 ;
        RECT 93.180 -12.330 94.710 -12.120 ;
        RECT 95.090 -12.210 95.540 -12.120 ;
        RECT 95.920 -12.330 97.450 -12.120 ;
        RECT 77.510 -12.780 77.960 -12.700 ;
        RECT 75.660 -13.020 77.960 -12.780 ;
        RECT 75.660 -13.120 76.110 -13.020 ;
        RECT 77.510 -13.120 77.960 -13.020 ;
        RECT 78.910 -12.780 79.360 -12.670 ;
        RECT 80.760 -12.780 81.210 -12.670 ;
        RECT 78.910 -13.020 81.210 -12.780 ;
        RECT 78.910 -13.090 79.360 -13.020 ;
        RECT 62.160 -13.650 62.610 -13.600 ;
        RECT 60.520 -13.940 62.610 -13.650 ;
        RECT 60.520 -13.990 60.970 -13.940 ;
        RECT 43.770 -14.570 44.220 -14.500 ;
        RECT 41.920 -14.810 44.220 -14.570 ;
        RECT 41.920 -14.920 42.370 -14.810 ;
        RECT 43.770 -14.920 44.220 -14.810 ;
        RECT 45.170 -14.570 45.620 -14.470 ;
        RECT 47.020 -14.570 47.470 -14.470 ;
        RECT 45.170 -14.810 47.470 -14.570 ;
        RECT 45.170 -14.890 45.620 -14.810 ;
        RECT 25.680 -15.470 27.210 -15.260 ;
        RECT 27.590 -15.470 28.040 -15.380 ;
        RECT 28.420 -15.470 29.950 -15.260 ;
        RECT 39.180 -15.260 39.630 -14.980 ;
        RECT 43.000 -15.260 43.450 -14.980 ;
        RECT 46.220 -15.250 46.630 -14.810 ;
        RECT 47.020 -14.920 47.470 -14.810 ;
        RECT 48.660 -14.570 49.110 -14.470 ;
        RECT 50.510 -14.570 50.960 -14.470 ;
        RECT 48.660 -14.810 50.960 -14.570 ;
        RECT 48.660 -14.920 49.110 -14.810 ;
        RECT 49.500 -15.250 49.910 -14.810 ;
        RECT 50.510 -14.890 50.960 -14.810 ;
        RECT 51.910 -14.570 52.360 -14.500 ;
        RECT 52.960 -14.570 53.370 -14.140 ;
        RECT 53.760 -14.570 54.210 -14.470 ;
        RECT 51.910 -14.810 54.210 -14.570 ;
        RECT 51.910 -14.920 52.360 -14.810 ;
        RECT 53.760 -14.920 54.210 -14.810 ;
        RECT 55.420 -14.570 55.870 -14.470 ;
        RECT 56.260 -14.570 56.670 -14.140 ;
        RECT 59.420 -14.210 60.970 -13.990 ;
        RECT 61.350 -14.000 61.780 -13.940 ;
        RECT 62.160 -13.990 62.610 -13.940 ;
        RECT 63.210 -13.990 63.710 -13.600 ;
        RECT 62.160 -14.210 63.710 -13.990 ;
        RECT 72.920 -13.600 74.470 -13.380 ;
        RECT 72.920 -13.990 73.420 -13.600 ;
        RECT 74.020 -13.650 74.470 -13.600 ;
        RECT 74.850 -13.650 75.280 -13.590 ;
        RECT 75.660 -13.600 77.210 -13.380 ;
        RECT 79.960 -13.450 80.370 -13.020 ;
        RECT 80.760 -13.120 81.210 -13.020 ;
        RECT 82.420 -12.780 82.870 -12.670 ;
        RECT 84.270 -12.780 84.720 -12.670 ;
        RECT 82.420 -13.020 84.720 -12.780 ;
        RECT 82.420 -13.120 82.870 -13.020 ;
        RECT 83.260 -13.450 83.670 -13.020 ;
        RECT 84.270 -13.090 84.720 -13.020 ;
        RECT 85.670 -12.780 86.120 -12.700 ;
        RECT 86.720 -12.780 87.130 -12.340 ;
        RECT 87.520 -12.780 87.970 -12.670 ;
        RECT 85.670 -13.020 87.970 -12.780 ;
        RECT 85.670 -13.120 86.120 -13.020 ;
        RECT 87.520 -13.120 87.970 -13.020 ;
        RECT 89.160 -12.780 89.610 -12.670 ;
        RECT 90.000 -12.780 90.410 -12.340 ;
        RECT 93.180 -12.610 93.630 -12.330 ;
        RECT 97.000 -12.610 97.450 -12.330 ;
        RECT 106.680 -12.170 110.950 -12.120 ;
        RECT 106.680 -12.330 108.210 -12.170 ;
        RECT 108.590 -12.210 109.040 -12.170 ;
        RECT 109.420 -12.330 110.950 -12.170 ;
        RECT 91.010 -12.780 91.460 -12.700 ;
        RECT 89.160 -13.020 91.460 -12.780 ;
        RECT 89.160 -13.120 89.610 -13.020 ;
        RECT 91.010 -13.120 91.460 -13.020 ;
        RECT 92.410 -12.780 92.860 -12.670 ;
        RECT 94.260 -12.780 94.710 -12.670 ;
        RECT 92.410 -13.020 94.710 -12.780 ;
        RECT 92.410 -13.090 92.860 -13.020 ;
        RECT 75.660 -13.650 76.110 -13.600 ;
        RECT 74.020 -13.940 76.110 -13.650 ;
        RECT 74.020 -13.990 74.470 -13.940 ;
        RECT 57.270 -14.570 57.720 -14.500 ;
        RECT 55.420 -14.810 57.720 -14.570 ;
        RECT 55.420 -14.920 55.870 -14.810 ;
        RECT 57.270 -14.920 57.720 -14.810 ;
        RECT 58.670 -14.570 59.120 -14.470 ;
        RECT 60.520 -14.570 60.970 -14.470 ;
        RECT 58.670 -14.810 60.970 -14.570 ;
        RECT 58.670 -14.890 59.120 -14.810 ;
        RECT 39.180 -15.470 40.710 -15.260 ;
        RECT 41.090 -15.470 41.540 -15.380 ;
        RECT 41.920 -15.470 43.450 -15.260 ;
        RECT 52.680 -15.260 53.130 -14.980 ;
        RECT 56.500 -15.260 56.950 -14.980 ;
        RECT 59.720 -15.250 60.130 -14.810 ;
        RECT 60.520 -14.920 60.970 -14.810 ;
        RECT 62.160 -14.570 62.610 -14.470 ;
        RECT 64.010 -14.570 64.460 -14.470 ;
        RECT 62.160 -14.810 64.460 -14.570 ;
        RECT 62.160 -14.920 62.610 -14.810 ;
        RECT 63.000 -15.250 63.410 -14.810 ;
        RECT 64.010 -14.890 64.460 -14.810 ;
        RECT 65.410 -14.570 65.860 -14.500 ;
        RECT 66.460 -14.570 66.870 -14.140 ;
        RECT 67.260 -14.570 67.710 -14.470 ;
        RECT 65.410 -14.810 67.710 -14.570 ;
        RECT 65.410 -14.920 65.860 -14.810 ;
        RECT 67.260 -14.920 67.710 -14.810 ;
        RECT 68.920 -14.570 69.370 -14.470 ;
        RECT 69.760 -14.570 70.170 -14.140 ;
        RECT 72.920 -14.210 74.470 -13.990 ;
        RECT 74.850 -14.000 75.280 -13.940 ;
        RECT 75.660 -13.990 76.110 -13.940 ;
        RECT 76.710 -13.990 77.210 -13.600 ;
        RECT 75.660 -14.210 77.210 -13.990 ;
        RECT 86.420 -13.600 87.970 -13.380 ;
        RECT 86.420 -13.990 86.920 -13.600 ;
        RECT 87.520 -13.650 87.970 -13.600 ;
        RECT 88.350 -13.650 88.780 -13.590 ;
        RECT 89.160 -13.600 90.710 -13.380 ;
        RECT 93.460 -13.450 93.870 -13.020 ;
        RECT 94.260 -13.120 94.710 -13.020 ;
        RECT 95.920 -12.780 96.370 -12.670 ;
        RECT 97.770 -12.780 98.220 -12.670 ;
        RECT 95.920 -13.020 98.220 -12.780 ;
        RECT 95.920 -13.120 96.370 -13.020 ;
        RECT 96.760 -13.450 97.170 -13.020 ;
        RECT 97.770 -13.090 98.220 -13.020 ;
        RECT 99.170 -12.780 99.620 -12.700 ;
        RECT 100.220 -12.780 100.630 -12.340 ;
        RECT 101.020 -12.780 101.470 -12.670 ;
        RECT 99.170 -13.020 101.470 -12.780 ;
        RECT 99.170 -13.120 99.620 -13.020 ;
        RECT 101.020 -13.120 101.470 -13.020 ;
        RECT 102.660 -12.780 103.110 -12.670 ;
        RECT 103.500 -12.780 103.910 -12.340 ;
        RECT 106.680 -12.610 107.130 -12.330 ;
        RECT 110.500 -12.610 110.950 -12.330 ;
        RECT 120.180 -12.330 121.710 -12.120 ;
        RECT 122.090 -12.210 122.540 -12.120 ;
        RECT 122.920 -12.330 124.450 -12.120 ;
        RECT 104.510 -12.780 104.960 -12.700 ;
        RECT 102.660 -13.020 104.960 -12.780 ;
        RECT 102.660 -13.120 103.110 -13.020 ;
        RECT 104.510 -13.120 104.960 -13.020 ;
        RECT 105.910 -12.780 106.360 -12.670 ;
        RECT 107.760 -12.780 108.210 -12.670 ;
        RECT 105.910 -13.020 108.210 -12.780 ;
        RECT 105.910 -13.090 106.360 -13.020 ;
        RECT 89.160 -13.650 89.610 -13.600 ;
        RECT 87.520 -13.940 89.610 -13.650 ;
        RECT 87.520 -13.990 87.970 -13.940 ;
        RECT 70.770 -14.570 71.220 -14.500 ;
        RECT 68.920 -14.810 71.220 -14.570 ;
        RECT 68.920 -14.920 69.370 -14.810 ;
        RECT 70.770 -14.920 71.220 -14.810 ;
        RECT 72.170 -14.570 72.620 -14.470 ;
        RECT 74.020 -14.570 74.470 -14.470 ;
        RECT 72.170 -14.810 74.470 -14.570 ;
        RECT 72.170 -14.890 72.620 -14.810 ;
        RECT 52.680 -15.470 54.210 -15.260 ;
        RECT 54.590 -15.470 55.040 -15.380 ;
        RECT 55.420 -15.470 56.950 -15.260 ;
        RECT 66.180 -15.260 66.630 -14.980 ;
        RECT 70.000 -15.260 70.450 -14.980 ;
        RECT 73.220 -15.250 73.630 -14.810 ;
        RECT 74.020 -14.920 74.470 -14.810 ;
        RECT 75.660 -14.570 76.110 -14.470 ;
        RECT 77.510 -14.570 77.960 -14.470 ;
        RECT 75.660 -14.810 77.960 -14.570 ;
        RECT 75.660 -14.920 76.110 -14.810 ;
        RECT 76.500 -15.250 76.910 -14.810 ;
        RECT 77.510 -14.890 77.960 -14.810 ;
        RECT 78.910 -14.570 79.360 -14.500 ;
        RECT 79.960 -14.570 80.370 -14.140 ;
        RECT 80.760 -14.570 81.210 -14.470 ;
        RECT 78.910 -14.810 81.210 -14.570 ;
        RECT 78.910 -14.920 79.360 -14.810 ;
        RECT 80.760 -14.920 81.210 -14.810 ;
        RECT 82.420 -14.570 82.870 -14.470 ;
        RECT 83.260 -14.570 83.670 -14.140 ;
        RECT 86.420 -14.210 87.970 -13.990 ;
        RECT 88.350 -14.000 88.780 -13.940 ;
        RECT 89.160 -13.990 89.610 -13.940 ;
        RECT 90.210 -13.990 90.710 -13.600 ;
        RECT 89.160 -14.210 90.710 -13.990 ;
        RECT 99.920 -13.600 101.470 -13.380 ;
        RECT 99.920 -13.990 100.420 -13.600 ;
        RECT 101.020 -13.650 101.470 -13.600 ;
        RECT 101.850 -13.650 102.280 -13.590 ;
        RECT 102.660 -13.600 104.210 -13.380 ;
        RECT 106.960 -13.450 107.370 -13.020 ;
        RECT 107.760 -13.120 108.210 -13.020 ;
        RECT 109.420 -12.780 109.870 -12.670 ;
        RECT 111.270 -12.780 111.720 -12.670 ;
        RECT 109.420 -13.020 111.720 -12.780 ;
        RECT 109.420 -13.120 109.870 -13.020 ;
        RECT 110.260 -13.450 110.670 -13.020 ;
        RECT 111.270 -13.090 111.720 -13.020 ;
        RECT 112.670 -12.780 113.120 -12.700 ;
        RECT 113.720 -12.780 114.130 -12.340 ;
        RECT 114.520 -12.780 114.970 -12.670 ;
        RECT 112.670 -13.020 114.970 -12.780 ;
        RECT 112.670 -13.120 113.120 -13.020 ;
        RECT 114.520 -13.120 114.970 -13.020 ;
        RECT 116.160 -12.780 116.610 -12.670 ;
        RECT 117.000 -12.780 117.410 -12.340 ;
        RECT 120.180 -12.610 120.630 -12.330 ;
        RECT 124.000 -12.610 124.450 -12.330 ;
        RECT 133.680 -12.330 135.210 -12.120 ;
        RECT 135.590 -12.210 136.040 -12.120 ;
        RECT 136.420 -12.330 137.950 -12.120 ;
        RECT 118.010 -12.780 118.460 -12.700 ;
        RECT 116.160 -13.020 118.460 -12.780 ;
        RECT 116.160 -13.120 116.610 -13.020 ;
        RECT 118.010 -13.120 118.460 -13.020 ;
        RECT 119.410 -12.780 119.860 -12.670 ;
        RECT 121.260 -12.780 121.710 -12.670 ;
        RECT 119.410 -13.020 121.710 -12.780 ;
        RECT 119.410 -13.090 119.860 -13.020 ;
        RECT 102.660 -13.650 103.110 -13.600 ;
        RECT 101.020 -13.940 103.110 -13.650 ;
        RECT 101.020 -13.990 101.470 -13.940 ;
        RECT 84.270 -14.570 84.720 -14.500 ;
        RECT 82.420 -14.810 84.720 -14.570 ;
        RECT 82.420 -14.920 82.870 -14.810 ;
        RECT 84.270 -14.920 84.720 -14.810 ;
        RECT 85.670 -14.570 86.120 -14.470 ;
        RECT 87.520 -14.570 87.970 -14.470 ;
        RECT 85.670 -14.810 87.970 -14.570 ;
        RECT 85.670 -14.890 86.120 -14.810 ;
        RECT 66.180 -15.470 67.710 -15.260 ;
        RECT 68.090 -15.470 68.540 -15.380 ;
        RECT 68.920 -15.470 70.450 -15.260 ;
        RECT 79.680 -15.260 80.130 -14.980 ;
        RECT 83.500 -15.260 83.950 -14.980 ;
        RECT 86.720 -15.250 87.130 -14.810 ;
        RECT 87.520 -14.920 87.970 -14.810 ;
        RECT 89.160 -14.570 89.610 -14.470 ;
        RECT 91.010 -14.570 91.460 -14.470 ;
        RECT 89.160 -14.810 91.460 -14.570 ;
        RECT 89.160 -14.920 89.610 -14.810 ;
        RECT 90.000 -15.250 90.410 -14.810 ;
        RECT 91.010 -14.890 91.460 -14.810 ;
        RECT 92.410 -14.570 92.860 -14.500 ;
        RECT 93.460 -14.570 93.870 -14.140 ;
        RECT 94.260 -14.570 94.710 -14.470 ;
        RECT 92.410 -14.810 94.710 -14.570 ;
        RECT 92.410 -14.920 92.860 -14.810 ;
        RECT 94.260 -14.920 94.710 -14.810 ;
        RECT 95.920 -14.570 96.370 -14.470 ;
        RECT 96.760 -14.570 97.170 -14.140 ;
        RECT 99.920 -14.210 101.470 -13.990 ;
        RECT 101.850 -14.000 102.280 -13.940 ;
        RECT 102.660 -13.990 103.110 -13.940 ;
        RECT 103.710 -13.990 104.210 -13.600 ;
        RECT 102.660 -14.210 104.210 -13.990 ;
        RECT 113.420 -13.600 114.970 -13.380 ;
        RECT 113.420 -13.990 113.920 -13.600 ;
        RECT 114.520 -13.650 114.970 -13.600 ;
        RECT 115.350 -13.650 115.780 -13.590 ;
        RECT 116.160 -13.600 117.710 -13.380 ;
        RECT 120.460 -13.450 120.870 -13.020 ;
        RECT 121.260 -13.120 121.710 -13.020 ;
        RECT 122.920 -12.780 123.370 -12.670 ;
        RECT 124.770 -12.780 125.220 -12.670 ;
        RECT 122.920 -13.020 125.220 -12.780 ;
        RECT 122.920 -13.120 123.370 -13.020 ;
        RECT 123.760 -13.450 124.170 -13.020 ;
        RECT 124.770 -13.090 125.220 -13.020 ;
        RECT 126.170 -12.780 126.620 -12.700 ;
        RECT 127.220 -12.780 127.630 -12.340 ;
        RECT 128.020 -12.780 128.470 -12.670 ;
        RECT 126.170 -13.020 128.470 -12.780 ;
        RECT 126.170 -13.120 126.620 -13.020 ;
        RECT 128.020 -13.120 128.470 -13.020 ;
        RECT 129.660 -12.780 130.110 -12.670 ;
        RECT 130.500 -12.780 130.910 -12.340 ;
        RECT 133.680 -12.610 134.130 -12.330 ;
        RECT 137.500 -12.610 137.950 -12.330 ;
        RECT 147.180 -12.330 148.710 -12.120 ;
        RECT 149.090 -12.210 149.540 -12.120 ;
        RECT 149.920 -12.330 151.450 -12.120 ;
        RECT 131.510 -12.780 131.960 -12.700 ;
        RECT 129.660 -13.020 131.960 -12.780 ;
        RECT 129.660 -13.120 130.110 -13.020 ;
        RECT 131.510 -13.120 131.960 -13.020 ;
        RECT 132.910 -12.780 133.360 -12.670 ;
        RECT 134.760 -12.780 135.210 -12.670 ;
        RECT 132.910 -13.020 135.210 -12.780 ;
        RECT 132.910 -13.090 133.360 -13.020 ;
        RECT 116.160 -13.650 116.610 -13.600 ;
        RECT 114.520 -13.940 116.610 -13.650 ;
        RECT 114.520 -13.990 114.970 -13.940 ;
        RECT 97.770 -14.570 98.220 -14.500 ;
        RECT 95.920 -14.810 98.220 -14.570 ;
        RECT 95.920 -14.920 96.370 -14.810 ;
        RECT 97.770 -14.920 98.220 -14.810 ;
        RECT 99.170 -14.570 99.620 -14.470 ;
        RECT 101.020 -14.570 101.470 -14.470 ;
        RECT 99.170 -14.810 101.470 -14.570 ;
        RECT 99.170 -14.890 99.620 -14.810 ;
        RECT 79.680 -15.470 81.210 -15.260 ;
        RECT 81.590 -15.470 82.040 -15.380 ;
        RECT 82.420 -15.470 83.950 -15.260 ;
        RECT 93.180 -15.260 93.630 -14.980 ;
        RECT 97.000 -15.260 97.450 -14.980 ;
        RECT 100.220 -15.250 100.630 -14.810 ;
        RECT 101.020 -14.920 101.470 -14.810 ;
        RECT 102.660 -14.570 103.110 -14.470 ;
        RECT 104.510 -14.570 104.960 -14.470 ;
        RECT 102.660 -14.810 104.960 -14.570 ;
        RECT 102.660 -14.920 103.110 -14.810 ;
        RECT 103.500 -15.250 103.910 -14.810 ;
        RECT 104.510 -14.890 104.960 -14.810 ;
        RECT 105.910 -14.570 106.360 -14.500 ;
        RECT 106.960 -14.570 107.370 -14.140 ;
        RECT 107.760 -14.570 108.210 -14.470 ;
        RECT 105.910 -14.810 108.210 -14.570 ;
        RECT 105.910 -14.920 106.360 -14.810 ;
        RECT 107.760 -14.920 108.210 -14.810 ;
        RECT 109.420 -14.570 109.870 -14.470 ;
        RECT 110.260 -14.570 110.670 -14.140 ;
        RECT 113.420 -14.210 114.970 -13.990 ;
        RECT 115.350 -14.000 115.780 -13.940 ;
        RECT 116.160 -13.990 116.610 -13.940 ;
        RECT 117.210 -13.990 117.710 -13.600 ;
        RECT 116.160 -14.210 117.710 -13.990 ;
        RECT 126.920 -13.600 128.470 -13.380 ;
        RECT 126.920 -13.990 127.420 -13.600 ;
        RECT 128.020 -13.650 128.470 -13.600 ;
        RECT 128.850 -13.650 129.280 -13.590 ;
        RECT 129.660 -13.600 131.210 -13.380 ;
        RECT 133.960 -13.450 134.370 -13.020 ;
        RECT 134.760 -13.120 135.210 -13.020 ;
        RECT 136.420 -12.780 136.870 -12.670 ;
        RECT 138.270 -12.780 138.720 -12.670 ;
        RECT 136.420 -13.020 138.720 -12.780 ;
        RECT 136.420 -13.120 136.870 -13.020 ;
        RECT 137.260 -13.450 137.670 -13.020 ;
        RECT 138.270 -13.090 138.720 -13.020 ;
        RECT 139.670 -12.780 140.120 -12.700 ;
        RECT 140.720 -12.780 141.130 -12.340 ;
        RECT 141.520 -12.780 141.970 -12.670 ;
        RECT 139.670 -13.020 141.970 -12.780 ;
        RECT 139.670 -13.120 140.120 -13.020 ;
        RECT 141.520 -13.120 141.970 -13.020 ;
        RECT 143.160 -12.780 143.610 -12.670 ;
        RECT 144.000 -12.780 144.410 -12.340 ;
        RECT 147.180 -12.610 147.630 -12.330 ;
        RECT 151.000 -12.610 151.450 -12.330 ;
        RECT 160.680 -12.170 164.950 -12.120 ;
        RECT 160.680 -12.330 162.210 -12.170 ;
        RECT 162.590 -12.210 163.040 -12.170 ;
        RECT 163.420 -12.330 164.950 -12.170 ;
        RECT 145.010 -12.780 145.460 -12.700 ;
        RECT 143.160 -13.020 145.460 -12.780 ;
        RECT 143.160 -13.120 143.610 -13.020 ;
        RECT 145.010 -13.120 145.460 -13.020 ;
        RECT 146.410 -12.780 146.860 -12.670 ;
        RECT 148.260 -12.780 148.710 -12.670 ;
        RECT 146.410 -13.020 148.710 -12.780 ;
        RECT 146.410 -13.090 146.860 -13.020 ;
        RECT 129.660 -13.650 130.110 -13.600 ;
        RECT 128.020 -13.940 130.110 -13.650 ;
        RECT 128.020 -13.990 128.470 -13.940 ;
        RECT 111.270 -14.570 111.720 -14.500 ;
        RECT 109.420 -14.810 111.720 -14.570 ;
        RECT 109.420 -14.920 109.870 -14.810 ;
        RECT 111.270 -14.920 111.720 -14.810 ;
        RECT 112.670 -14.570 113.120 -14.470 ;
        RECT 114.520 -14.570 114.970 -14.470 ;
        RECT 112.670 -14.810 114.970 -14.570 ;
        RECT 112.670 -14.890 113.120 -14.810 ;
        RECT 93.180 -15.470 94.710 -15.260 ;
        RECT 95.090 -15.470 95.540 -15.380 ;
        RECT 95.920 -15.470 97.450 -15.260 ;
        RECT 106.680 -15.260 107.130 -14.980 ;
        RECT 110.500 -15.260 110.950 -14.980 ;
        RECT 113.720 -15.250 114.130 -14.810 ;
        RECT 114.520 -14.920 114.970 -14.810 ;
        RECT 116.160 -14.570 116.610 -14.470 ;
        RECT 118.010 -14.570 118.460 -14.470 ;
        RECT 116.160 -14.810 118.460 -14.570 ;
        RECT 116.160 -14.920 116.610 -14.810 ;
        RECT 117.000 -15.250 117.410 -14.810 ;
        RECT 118.010 -14.890 118.460 -14.810 ;
        RECT 119.410 -14.570 119.860 -14.500 ;
        RECT 120.460 -14.570 120.870 -14.140 ;
        RECT 121.260 -14.570 121.710 -14.470 ;
        RECT 119.410 -14.810 121.710 -14.570 ;
        RECT 119.410 -14.920 119.860 -14.810 ;
        RECT 121.260 -14.920 121.710 -14.810 ;
        RECT 122.920 -14.570 123.370 -14.470 ;
        RECT 123.760 -14.570 124.170 -14.140 ;
        RECT 126.920 -14.210 128.470 -13.990 ;
        RECT 128.850 -14.000 129.280 -13.940 ;
        RECT 129.660 -13.990 130.110 -13.940 ;
        RECT 130.710 -13.990 131.210 -13.600 ;
        RECT 129.660 -14.210 131.210 -13.990 ;
        RECT 140.420 -13.600 141.970 -13.380 ;
        RECT 140.420 -13.990 140.920 -13.600 ;
        RECT 141.520 -13.650 141.970 -13.600 ;
        RECT 142.350 -13.650 142.780 -13.590 ;
        RECT 143.160 -13.600 144.710 -13.380 ;
        RECT 147.460 -13.450 147.870 -13.020 ;
        RECT 148.260 -13.120 148.710 -13.020 ;
        RECT 149.920 -12.780 150.370 -12.670 ;
        RECT 151.770 -12.780 152.220 -12.670 ;
        RECT 149.920 -13.020 152.220 -12.780 ;
        RECT 149.920 -13.120 150.370 -13.020 ;
        RECT 150.760 -13.450 151.170 -13.020 ;
        RECT 151.770 -13.090 152.220 -13.020 ;
        RECT 153.170 -12.780 153.620 -12.700 ;
        RECT 154.220 -12.780 154.630 -12.340 ;
        RECT 155.020 -12.780 155.470 -12.670 ;
        RECT 153.170 -13.020 155.470 -12.780 ;
        RECT 153.170 -13.120 153.620 -13.020 ;
        RECT 155.020 -13.120 155.470 -13.020 ;
        RECT 156.660 -12.780 157.110 -12.670 ;
        RECT 157.500 -12.780 157.910 -12.340 ;
        RECT 160.680 -12.610 161.130 -12.330 ;
        RECT 164.500 -12.610 164.950 -12.330 ;
        RECT 174.180 -12.330 175.710 -12.120 ;
        RECT 176.090 -12.210 176.540 -12.120 ;
        RECT 176.920 -12.330 178.450 -12.120 ;
        RECT 158.510 -12.780 158.960 -12.700 ;
        RECT 156.660 -13.020 158.960 -12.780 ;
        RECT 156.660 -13.120 157.110 -13.020 ;
        RECT 158.510 -13.120 158.960 -13.020 ;
        RECT 159.910 -12.780 160.360 -12.670 ;
        RECT 161.760 -12.780 162.210 -12.670 ;
        RECT 159.910 -13.020 162.210 -12.780 ;
        RECT 159.910 -13.090 160.360 -13.020 ;
        RECT 143.160 -13.650 143.610 -13.600 ;
        RECT 141.520 -13.940 143.610 -13.650 ;
        RECT 141.520 -13.990 141.970 -13.940 ;
        RECT 124.770 -14.570 125.220 -14.500 ;
        RECT 122.920 -14.810 125.220 -14.570 ;
        RECT 122.920 -14.920 123.370 -14.810 ;
        RECT 124.770 -14.920 125.220 -14.810 ;
        RECT 126.170 -14.570 126.620 -14.470 ;
        RECT 128.020 -14.570 128.470 -14.470 ;
        RECT 126.170 -14.810 128.470 -14.570 ;
        RECT 126.170 -14.890 126.620 -14.810 ;
        RECT 106.680 -15.470 108.210 -15.260 ;
        RECT 108.590 -15.470 109.040 -15.380 ;
        RECT 109.420 -15.470 110.950 -15.260 ;
        RECT 120.180 -15.260 120.630 -14.980 ;
        RECT 124.000 -15.260 124.450 -14.980 ;
        RECT 127.220 -15.250 127.630 -14.810 ;
        RECT 128.020 -14.920 128.470 -14.810 ;
        RECT 129.660 -14.570 130.110 -14.470 ;
        RECT 131.510 -14.570 131.960 -14.470 ;
        RECT 129.660 -14.810 131.960 -14.570 ;
        RECT 129.660 -14.920 130.110 -14.810 ;
        RECT 130.500 -15.250 130.910 -14.810 ;
        RECT 131.510 -14.890 131.960 -14.810 ;
        RECT 132.910 -14.570 133.360 -14.500 ;
        RECT 133.960 -14.570 134.370 -14.140 ;
        RECT 134.760 -14.570 135.210 -14.470 ;
        RECT 132.910 -14.810 135.210 -14.570 ;
        RECT 132.910 -14.920 133.360 -14.810 ;
        RECT 134.760 -14.920 135.210 -14.810 ;
        RECT 136.420 -14.570 136.870 -14.470 ;
        RECT 137.260 -14.570 137.670 -14.140 ;
        RECT 140.420 -14.210 141.970 -13.990 ;
        RECT 142.350 -14.000 142.780 -13.940 ;
        RECT 143.160 -13.990 143.610 -13.940 ;
        RECT 144.210 -13.990 144.710 -13.600 ;
        RECT 143.160 -14.210 144.710 -13.990 ;
        RECT 153.920 -13.600 155.470 -13.380 ;
        RECT 153.920 -13.990 154.420 -13.600 ;
        RECT 155.020 -13.650 155.470 -13.600 ;
        RECT 155.850 -13.650 156.280 -13.590 ;
        RECT 156.660 -13.600 158.210 -13.380 ;
        RECT 160.960 -13.450 161.370 -13.020 ;
        RECT 161.760 -13.120 162.210 -13.020 ;
        RECT 163.420 -12.780 163.870 -12.670 ;
        RECT 165.270 -12.780 165.720 -12.670 ;
        RECT 163.420 -13.020 165.720 -12.780 ;
        RECT 163.420 -13.120 163.870 -13.020 ;
        RECT 164.260 -13.450 164.670 -13.020 ;
        RECT 165.270 -13.090 165.720 -13.020 ;
        RECT 166.670 -12.780 167.120 -12.700 ;
        RECT 167.720 -12.780 168.130 -12.340 ;
        RECT 168.520 -12.780 168.970 -12.670 ;
        RECT 166.670 -13.020 168.970 -12.780 ;
        RECT 166.670 -13.120 167.120 -13.020 ;
        RECT 168.520 -13.120 168.970 -13.020 ;
        RECT 170.160 -12.780 170.610 -12.670 ;
        RECT 171.000 -12.780 171.410 -12.340 ;
        RECT 174.180 -12.610 174.630 -12.330 ;
        RECT 178.000 -12.610 178.450 -12.330 ;
        RECT 187.680 -12.330 189.210 -12.120 ;
        RECT 189.590 -12.210 190.040 -12.120 ;
        RECT 190.420 -12.330 191.950 -12.120 ;
        RECT 172.010 -12.780 172.460 -12.700 ;
        RECT 170.160 -13.020 172.460 -12.780 ;
        RECT 170.160 -13.120 170.610 -13.020 ;
        RECT 172.010 -13.120 172.460 -13.020 ;
        RECT 173.410 -12.780 173.860 -12.670 ;
        RECT 175.260 -12.780 175.710 -12.670 ;
        RECT 173.410 -13.020 175.710 -12.780 ;
        RECT 173.410 -13.090 173.860 -13.020 ;
        RECT 156.660 -13.650 157.110 -13.600 ;
        RECT 155.020 -13.940 157.110 -13.650 ;
        RECT 155.020 -13.990 155.470 -13.940 ;
        RECT 138.270 -14.570 138.720 -14.500 ;
        RECT 136.420 -14.810 138.720 -14.570 ;
        RECT 136.420 -14.920 136.870 -14.810 ;
        RECT 138.270 -14.920 138.720 -14.810 ;
        RECT 139.670 -14.570 140.120 -14.470 ;
        RECT 141.520 -14.570 141.970 -14.470 ;
        RECT 139.670 -14.810 141.970 -14.570 ;
        RECT 139.670 -14.890 140.120 -14.810 ;
        RECT 120.180 -15.470 121.710 -15.260 ;
        RECT 122.090 -15.470 122.540 -15.380 ;
        RECT 122.920 -15.470 124.450 -15.260 ;
        RECT 133.680 -15.260 134.130 -14.980 ;
        RECT 137.500 -15.260 137.950 -14.980 ;
        RECT 140.720 -15.250 141.130 -14.810 ;
        RECT 141.520 -14.920 141.970 -14.810 ;
        RECT 143.160 -14.570 143.610 -14.470 ;
        RECT 145.010 -14.570 145.460 -14.470 ;
        RECT 143.160 -14.810 145.460 -14.570 ;
        RECT 143.160 -14.920 143.610 -14.810 ;
        RECT 144.000 -15.250 144.410 -14.810 ;
        RECT 145.010 -14.890 145.460 -14.810 ;
        RECT 146.410 -14.570 146.860 -14.500 ;
        RECT 147.460 -14.570 147.870 -14.140 ;
        RECT 148.260 -14.570 148.710 -14.470 ;
        RECT 146.410 -14.810 148.710 -14.570 ;
        RECT 146.410 -14.920 146.860 -14.810 ;
        RECT 148.260 -14.920 148.710 -14.810 ;
        RECT 149.920 -14.570 150.370 -14.470 ;
        RECT 150.760 -14.570 151.170 -14.140 ;
        RECT 153.920 -14.210 155.470 -13.990 ;
        RECT 155.850 -14.000 156.280 -13.940 ;
        RECT 156.660 -13.990 157.110 -13.940 ;
        RECT 157.710 -13.990 158.210 -13.600 ;
        RECT 156.660 -14.210 158.210 -13.990 ;
        RECT 167.420 -13.600 168.970 -13.380 ;
        RECT 167.420 -13.990 167.920 -13.600 ;
        RECT 168.520 -13.650 168.970 -13.600 ;
        RECT 169.350 -13.650 169.780 -13.590 ;
        RECT 170.160 -13.600 171.710 -13.380 ;
        RECT 174.460 -13.450 174.870 -13.020 ;
        RECT 175.260 -13.120 175.710 -13.020 ;
        RECT 176.920 -12.780 177.370 -12.670 ;
        RECT 178.770 -12.780 179.220 -12.670 ;
        RECT 176.920 -13.020 179.220 -12.780 ;
        RECT 176.920 -13.120 177.370 -13.020 ;
        RECT 177.760 -13.450 178.170 -13.020 ;
        RECT 178.770 -13.090 179.220 -13.020 ;
        RECT 180.170 -12.780 180.620 -12.700 ;
        RECT 181.220 -12.780 181.630 -12.340 ;
        RECT 182.020 -12.780 182.470 -12.670 ;
        RECT 180.170 -13.020 182.470 -12.780 ;
        RECT 180.170 -13.120 180.620 -13.020 ;
        RECT 182.020 -13.120 182.470 -13.020 ;
        RECT 183.660 -12.780 184.110 -12.670 ;
        RECT 184.500 -12.780 184.910 -12.340 ;
        RECT 187.680 -12.610 188.130 -12.330 ;
        RECT 191.500 -12.610 191.950 -12.330 ;
        RECT 201.180 -12.330 202.710 -12.120 ;
        RECT 203.090 -12.210 203.540 -12.120 ;
        RECT 203.920 -12.330 205.450 -12.120 ;
        RECT 185.510 -12.780 185.960 -12.700 ;
        RECT 183.660 -13.020 185.960 -12.780 ;
        RECT 183.660 -13.120 184.110 -13.020 ;
        RECT 185.510 -13.120 185.960 -13.020 ;
        RECT 186.910 -12.780 187.360 -12.670 ;
        RECT 188.760 -12.780 189.210 -12.670 ;
        RECT 186.910 -13.020 189.210 -12.780 ;
        RECT 186.910 -13.090 187.360 -13.020 ;
        RECT 170.160 -13.650 170.610 -13.600 ;
        RECT 168.520 -13.940 170.610 -13.650 ;
        RECT 168.520 -13.990 168.970 -13.940 ;
        RECT 151.770 -14.570 152.220 -14.500 ;
        RECT 149.920 -14.810 152.220 -14.570 ;
        RECT 149.920 -14.920 150.370 -14.810 ;
        RECT 151.770 -14.920 152.220 -14.810 ;
        RECT 153.170 -14.570 153.620 -14.470 ;
        RECT 155.020 -14.570 155.470 -14.470 ;
        RECT 153.170 -14.810 155.470 -14.570 ;
        RECT 153.170 -14.890 153.620 -14.810 ;
        RECT 133.680 -15.470 135.210 -15.260 ;
        RECT 135.590 -15.470 136.040 -15.380 ;
        RECT 136.420 -15.470 137.950 -15.260 ;
        RECT 147.180 -15.260 147.630 -14.980 ;
        RECT 151.000 -15.260 151.450 -14.980 ;
        RECT 154.220 -15.250 154.630 -14.810 ;
        RECT 155.020 -14.920 155.470 -14.810 ;
        RECT 156.660 -14.570 157.110 -14.470 ;
        RECT 158.510 -14.570 158.960 -14.470 ;
        RECT 156.660 -14.810 158.960 -14.570 ;
        RECT 156.660 -14.920 157.110 -14.810 ;
        RECT 157.500 -15.250 157.910 -14.810 ;
        RECT 158.510 -14.890 158.960 -14.810 ;
        RECT 159.910 -14.570 160.360 -14.500 ;
        RECT 160.960 -14.570 161.370 -14.140 ;
        RECT 161.760 -14.570 162.210 -14.470 ;
        RECT 159.910 -14.810 162.210 -14.570 ;
        RECT 159.910 -14.920 160.360 -14.810 ;
        RECT 161.760 -14.920 162.210 -14.810 ;
        RECT 163.420 -14.570 163.870 -14.470 ;
        RECT 164.260 -14.570 164.670 -14.140 ;
        RECT 167.420 -14.210 168.970 -13.990 ;
        RECT 169.350 -14.000 169.780 -13.940 ;
        RECT 170.160 -13.990 170.610 -13.940 ;
        RECT 171.210 -13.990 171.710 -13.600 ;
        RECT 170.160 -14.210 171.710 -13.990 ;
        RECT 180.920 -13.600 182.470 -13.380 ;
        RECT 180.920 -13.990 181.420 -13.600 ;
        RECT 182.020 -13.650 182.470 -13.600 ;
        RECT 182.850 -13.650 183.280 -13.590 ;
        RECT 183.660 -13.600 185.210 -13.380 ;
        RECT 187.960 -13.450 188.370 -13.020 ;
        RECT 188.760 -13.120 189.210 -13.020 ;
        RECT 190.420 -12.780 190.870 -12.670 ;
        RECT 192.270 -12.780 192.720 -12.670 ;
        RECT 190.420 -13.020 192.720 -12.780 ;
        RECT 190.420 -13.120 190.870 -13.020 ;
        RECT 191.260 -13.450 191.670 -13.020 ;
        RECT 192.270 -13.090 192.720 -13.020 ;
        RECT 193.670 -12.780 194.120 -12.700 ;
        RECT 194.720 -12.780 195.130 -12.340 ;
        RECT 195.520 -12.780 195.970 -12.670 ;
        RECT 193.670 -13.020 195.970 -12.780 ;
        RECT 193.670 -13.120 194.120 -13.020 ;
        RECT 195.520 -13.120 195.970 -13.020 ;
        RECT 197.160 -12.780 197.610 -12.670 ;
        RECT 198.000 -12.780 198.410 -12.340 ;
        RECT 201.180 -12.610 201.630 -12.330 ;
        RECT 205.000 -12.610 205.450 -12.330 ;
        RECT 214.680 -12.330 216.210 -12.120 ;
        RECT 216.590 -12.170 217.690 -12.120 ;
        RECT 216.590 -12.210 217.030 -12.170 ;
        RECT 199.010 -12.780 199.460 -12.700 ;
        RECT 197.160 -13.020 199.460 -12.780 ;
        RECT 197.160 -13.120 197.610 -13.020 ;
        RECT 199.010 -13.120 199.460 -13.020 ;
        RECT 200.410 -12.780 200.860 -12.670 ;
        RECT 202.260 -12.780 202.710 -12.670 ;
        RECT 200.410 -13.020 202.710 -12.780 ;
        RECT 200.410 -13.090 200.860 -13.020 ;
        RECT 183.660 -13.650 184.110 -13.600 ;
        RECT 182.020 -13.940 184.110 -13.650 ;
        RECT 182.020 -13.990 182.470 -13.940 ;
        RECT 165.270 -14.570 165.720 -14.500 ;
        RECT 163.420 -14.810 165.720 -14.570 ;
        RECT 163.420 -14.920 163.870 -14.810 ;
        RECT 165.270 -14.920 165.720 -14.810 ;
        RECT 166.670 -14.570 167.120 -14.470 ;
        RECT 168.520 -14.570 168.970 -14.470 ;
        RECT 166.670 -14.810 168.970 -14.570 ;
        RECT 166.670 -14.890 167.120 -14.810 ;
        RECT 147.180 -15.470 148.710 -15.260 ;
        RECT 149.090 -15.470 149.540 -15.380 ;
        RECT 149.920 -15.470 151.450 -15.260 ;
        RECT 160.680 -15.260 161.130 -14.980 ;
        RECT 164.500 -15.260 164.950 -14.980 ;
        RECT 167.720 -15.250 168.130 -14.810 ;
        RECT 168.520 -14.920 168.970 -14.810 ;
        RECT 170.160 -14.570 170.610 -14.470 ;
        RECT 172.010 -14.570 172.460 -14.470 ;
        RECT 170.160 -14.810 172.460 -14.570 ;
        RECT 170.160 -14.920 170.610 -14.810 ;
        RECT 171.000 -15.250 171.410 -14.810 ;
        RECT 172.010 -14.890 172.460 -14.810 ;
        RECT 173.410 -14.570 173.860 -14.500 ;
        RECT 174.460 -14.570 174.870 -14.140 ;
        RECT 175.260 -14.570 175.710 -14.470 ;
        RECT 173.410 -14.810 175.710 -14.570 ;
        RECT 173.410 -14.920 173.860 -14.810 ;
        RECT 175.260 -14.920 175.710 -14.810 ;
        RECT 176.920 -14.570 177.370 -14.470 ;
        RECT 177.760 -14.570 178.170 -14.140 ;
        RECT 180.920 -14.210 182.470 -13.990 ;
        RECT 182.850 -14.000 183.280 -13.940 ;
        RECT 183.660 -13.990 184.110 -13.940 ;
        RECT 184.710 -13.990 185.210 -13.600 ;
        RECT 183.660 -14.210 185.210 -13.990 ;
        RECT 194.420 -13.600 195.970 -13.380 ;
        RECT 194.420 -13.990 194.920 -13.600 ;
        RECT 195.520 -13.650 195.970 -13.600 ;
        RECT 196.350 -13.650 196.780 -13.590 ;
        RECT 197.160 -13.600 198.710 -13.380 ;
        RECT 201.460 -13.450 201.870 -13.020 ;
        RECT 202.260 -13.120 202.710 -13.020 ;
        RECT 203.920 -12.780 204.370 -12.670 ;
        RECT 205.770 -12.780 206.220 -12.670 ;
        RECT 203.920 -13.020 206.220 -12.780 ;
        RECT 203.920 -13.120 204.370 -13.020 ;
        RECT 204.760 -13.450 205.170 -13.020 ;
        RECT 205.770 -13.090 206.220 -13.020 ;
        RECT 207.170 -12.780 207.620 -12.700 ;
        RECT 208.220 -12.780 208.630 -12.340 ;
        RECT 209.020 -12.780 209.470 -12.670 ;
        RECT 207.170 -13.020 209.470 -12.780 ;
        RECT 207.170 -13.120 207.620 -13.020 ;
        RECT 209.020 -13.120 209.470 -13.020 ;
        RECT 210.660 -12.780 211.110 -12.670 ;
        RECT 211.500 -12.780 211.910 -12.340 ;
        RECT 214.680 -12.610 215.130 -12.330 ;
        RECT 212.510 -12.780 212.960 -12.700 ;
        RECT 210.660 -13.020 212.960 -12.780 ;
        RECT 210.660 -13.120 211.110 -13.020 ;
        RECT 212.510 -13.120 212.960 -13.020 ;
        RECT 213.910 -12.780 214.360 -12.670 ;
        RECT 215.760 -12.780 216.210 -12.670 ;
        RECT 213.910 -13.020 216.210 -12.780 ;
        RECT 213.910 -13.090 214.360 -13.020 ;
        RECT 197.160 -13.650 197.610 -13.600 ;
        RECT 195.520 -13.940 197.610 -13.650 ;
        RECT 195.520 -13.990 195.970 -13.940 ;
        RECT 178.770 -14.570 179.220 -14.500 ;
        RECT 176.920 -14.810 179.220 -14.570 ;
        RECT 176.920 -14.920 177.370 -14.810 ;
        RECT 178.770 -14.920 179.220 -14.810 ;
        RECT 180.170 -14.570 180.620 -14.470 ;
        RECT 182.020 -14.570 182.470 -14.470 ;
        RECT 180.170 -14.810 182.470 -14.570 ;
        RECT 180.170 -14.890 180.620 -14.810 ;
        RECT 160.680 -15.470 162.210 -15.260 ;
        RECT 162.590 -15.470 163.040 -15.380 ;
        RECT 163.420 -15.470 164.950 -15.260 ;
        RECT 174.180 -15.260 174.630 -14.980 ;
        RECT 178.000 -15.260 178.450 -14.980 ;
        RECT 181.220 -15.250 181.630 -14.810 ;
        RECT 182.020 -14.920 182.470 -14.810 ;
        RECT 183.660 -14.570 184.110 -14.470 ;
        RECT 185.510 -14.570 185.960 -14.470 ;
        RECT 183.660 -14.810 185.960 -14.570 ;
        RECT 183.660 -14.920 184.110 -14.810 ;
        RECT 184.500 -15.250 184.910 -14.810 ;
        RECT 185.510 -14.890 185.960 -14.810 ;
        RECT 186.910 -14.570 187.360 -14.500 ;
        RECT 187.960 -14.570 188.370 -14.140 ;
        RECT 188.760 -14.570 189.210 -14.470 ;
        RECT 186.910 -14.810 189.210 -14.570 ;
        RECT 186.910 -14.920 187.360 -14.810 ;
        RECT 188.760 -14.920 189.210 -14.810 ;
        RECT 190.420 -14.570 190.870 -14.470 ;
        RECT 191.260 -14.570 191.670 -14.140 ;
        RECT 194.420 -14.210 195.970 -13.990 ;
        RECT 196.350 -14.000 196.780 -13.940 ;
        RECT 197.160 -13.990 197.610 -13.940 ;
        RECT 198.210 -13.990 198.710 -13.600 ;
        RECT 197.160 -14.210 198.710 -13.990 ;
        RECT 207.920 -13.600 209.470 -13.380 ;
        RECT 207.920 -13.990 208.420 -13.600 ;
        RECT 209.020 -13.650 209.470 -13.600 ;
        RECT 209.850 -13.650 210.280 -13.590 ;
        RECT 210.660 -13.600 212.210 -13.380 ;
        RECT 214.960 -13.450 215.370 -13.020 ;
        RECT 215.760 -13.120 216.210 -13.020 ;
        RECT 210.660 -13.650 211.110 -13.600 ;
        RECT 209.020 -13.940 211.110 -13.650 ;
        RECT 209.020 -13.990 209.470 -13.940 ;
        RECT 192.270 -14.570 192.720 -14.500 ;
        RECT 190.420 -14.810 192.720 -14.570 ;
        RECT 190.420 -14.920 190.870 -14.810 ;
        RECT 192.270 -14.920 192.720 -14.810 ;
        RECT 193.670 -14.570 194.120 -14.470 ;
        RECT 195.520 -14.570 195.970 -14.470 ;
        RECT 193.670 -14.810 195.970 -14.570 ;
        RECT 193.670 -14.890 194.120 -14.810 ;
        RECT 174.180 -15.470 175.710 -15.260 ;
        RECT 176.090 -15.470 176.540 -15.380 ;
        RECT 176.920 -15.470 178.450 -15.260 ;
        RECT 187.680 -15.260 188.130 -14.980 ;
        RECT 191.500 -15.260 191.950 -14.980 ;
        RECT 194.720 -15.250 195.130 -14.810 ;
        RECT 195.520 -14.920 195.970 -14.810 ;
        RECT 197.160 -14.570 197.610 -14.470 ;
        RECT 199.010 -14.570 199.460 -14.470 ;
        RECT 197.160 -14.810 199.460 -14.570 ;
        RECT 197.160 -14.920 197.610 -14.810 ;
        RECT 198.000 -15.250 198.410 -14.810 ;
        RECT 199.010 -14.890 199.460 -14.810 ;
        RECT 200.410 -14.570 200.860 -14.500 ;
        RECT 201.460 -14.570 201.870 -14.140 ;
        RECT 202.260 -14.570 202.710 -14.470 ;
        RECT 200.410 -14.810 202.710 -14.570 ;
        RECT 200.410 -14.920 200.860 -14.810 ;
        RECT 202.260 -14.920 202.710 -14.810 ;
        RECT 203.920 -14.570 204.370 -14.470 ;
        RECT 204.760 -14.570 205.170 -14.140 ;
        RECT 207.920 -14.210 209.470 -13.990 ;
        RECT 209.850 -14.000 210.280 -13.940 ;
        RECT 210.660 -13.990 211.110 -13.940 ;
        RECT 211.710 -13.990 212.210 -13.600 ;
        RECT 210.660 -14.210 212.210 -13.990 ;
        RECT 205.770 -14.570 206.220 -14.500 ;
        RECT 203.920 -14.810 206.220 -14.570 ;
        RECT 203.920 -14.920 204.370 -14.810 ;
        RECT 205.770 -14.920 206.220 -14.810 ;
        RECT 207.170 -14.570 207.620 -14.470 ;
        RECT 209.020 -14.570 209.470 -14.470 ;
        RECT 207.170 -14.810 209.470 -14.570 ;
        RECT 207.170 -14.890 207.620 -14.810 ;
        RECT 187.680 -15.470 189.210 -15.260 ;
        RECT 189.590 -15.470 190.040 -15.380 ;
        RECT 190.420 -15.470 191.950 -15.260 ;
        RECT 201.180 -15.260 201.630 -14.980 ;
        RECT 205.000 -15.260 205.450 -14.980 ;
        RECT 208.220 -15.250 208.630 -14.810 ;
        RECT 209.020 -14.920 209.470 -14.810 ;
        RECT 210.660 -14.570 211.110 -14.470 ;
        RECT 212.510 -14.570 212.960 -14.470 ;
        RECT 210.660 -14.810 212.960 -14.570 ;
        RECT 210.660 -14.920 211.110 -14.810 ;
        RECT 211.500 -15.250 211.910 -14.810 ;
        RECT 212.510 -14.890 212.960 -14.810 ;
        RECT 213.910 -14.570 214.360 -14.500 ;
        RECT 214.960 -14.570 215.370 -14.140 ;
        RECT 215.760 -14.570 216.210 -14.470 ;
        RECT 213.910 -14.810 216.210 -14.570 ;
        RECT 213.910 -14.920 214.360 -14.810 ;
        RECT 215.760 -14.920 216.210 -14.810 ;
        RECT 201.180 -15.470 202.710 -15.260 ;
        RECT 203.090 -15.470 203.540 -15.380 ;
        RECT 203.920 -15.470 205.450 -15.260 ;
        RECT 214.680 -15.260 215.130 -14.980 ;
        RECT 214.680 -15.470 216.210 -15.260 ;
        RECT 216.590 -15.470 217.030 -15.380 ;
        RECT 13.260 -15.730 15.370 -15.470 ;
        RECT 26.760 -15.730 28.870 -15.470 ;
        RECT 40.260 -15.730 42.370 -15.470 ;
        RECT 53.760 -15.730 55.870 -15.470 ;
        RECT 67.260 -15.730 69.370 -15.470 ;
        RECT 80.760 -15.730 82.870 -15.470 ;
        RECT 94.260 -15.730 96.370 -15.470 ;
        RECT 107.760 -15.730 109.870 -15.470 ;
        RECT 121.260 -15.730 123.370 -15.470 ;
        RECT 134.760 -15.730 136.870 -15.470 ;
        RECT 148.260 -15.730 150.370 -15.470 ;
        RECT 161.760 -15.730 163.870 -15.470 ;
        RECT 175.260 -15.730 177.370 -15.470 ;
        RECT 188.760 -15.730 190.870 -15.470 ;
        RECT 202.260 -15.730 204.370 -15.470 ;
        RECT 215.760 -15.480 217.030 -15.470 ;
        RECT 215.760 -15.670 217.240 -15.480 ;
        RECT 215.760 -15.730 217.030 -15.670 ;
        RECT 12.180 -15.940 13.710 -15.730 ;
        RECT 14.090 -15.820 14.540 -15.730 ;
        RECT 14.920 -15.940 16.450 -15.730 ;
        RECT 1.420 -16.390 1.870 -16.280 ;
        RECT 3.270 -16.390 3.720 -16.280 ;
        RECT 1.420 -16.630 3.720 -16.390 ;
        RECT 1.420 -16.730 1.870 -16.630 ;
        RECT 2.260 -17.060 2.670 -16.630 ;
        RECT 3.270 -16.700 3.720 -16.630 ;
        RECT 4.670 -16.390 5.120 -16.310 ;
        RECT 5.720 -16.390 6.130 -15.950 ;
        RECT 6.520 -16.390 6.970 -16.280 ;
        RECT 4.670 -16.630 6.970 -16.390 ;
        RECT 4.670 -16.730 5.120 -16.630 ;
        RECT 6.520 -16.730 6.970 -16.630 ;
        RECT 8.160 -16.390 8.610 -16.280 ;
        RECT 9.000 -16.390 9.410 -15.950 ;
        RECT 12.180 -16.220 12.630 -15.940 ;
        RECT 16.000 -16.220 16.450 -15.940 ;
        RECT 25.680 -15.940 27.210 -15.730 ;
        RECT 27.590 -15.820 28.040 -15.730 ;
        RECT 28.420 -15.940 29.950 -15.730 ;
        RECT 10.010 -16.390 10.460 -16.310 ;
        RECT 8.160 -16.630 10.460 -16.390 ;
        RECT 8.160 -16.730 8.610 -16.630 ;
        RECT 10.010 -16.730 10.460 -16.630 ;
        RECT 11.410 -16.390 11.860 -16.280 ;
        RECT 13.260 -16.390 13.710 -16.280 ;
        RECT 11.410 -16.630 13.710 -16.390 ;
        RECT 11.410 -16.700 11.860 -16.630 ;
        RECT 5.420 -17.210 6.970 -16.990 ;
        RECT 5.420 -17.600 5.920 -17.210 ;
        RECT 6.520 -17.260 6.970 -17.210 ;
        RECT 7.350 -17.260 7.780 -17.200 ;
        RECT 8.160 -17.210 9.710 -16.990 ;
        RECT 12.460 -17.060 12.870 -16.630 ;
        RECT 13.260 -16.730 13.710 -16.630 ;
        RECT 14.920 -16.390 15.370 -16.280 ;
        RECT 16.770 -16.390 17.220 -16.280 ;
        RECT 14.920 -16.630 17.220 -16.390 ;
        RECT 14.920 -16.730 15.370 -16.630 ;
        RECT 15.760 -17.060 16.170 -16.630 ;
        RECT 16.770 -16.700 17.220 -16.630 ;
        RECT 18.170 -16.390 18.620 -16.310 ;
        RECT 19.220 -16.390 19.630 -15.950 ;
        RECT 20.020 -16.390 20.470 -16.280 ;
        RECT 18.170 -16.630 20.470 -16.390 ;
        RECT 18.170 -16.730 18.620 -16.630 ;
        RECT 20.020 -16.730 20.470 -16.630 ;
        RECT 21.660 -16.390 22.110 -16.280 ;
        RECT 22.500 -16.390 22.910 -15.950 ;
        RECT 25.680 -16.220 26.130 -15.940 ;
        RECT 29.500 -16.220 29.950 -15.940 ;
        RECT 39.180 -15.940 40.710 -15.730 ;
        RECT 41.090 -15.820 41.540 -15.730 ;
        RECT 41.920 -15.940 43.450 -15.730 ;
        RECT 23.510 -16.390 23.960 -16.310 ;
        RECT 21.660 -16.630 23.960 -16.390 ;
        RECT 21.660 -16.730 22.110 -16.630 ;
        RECT 23.510 -16.730 23.960 -16.630 ;
        RECT 24.910 -16.390 25.360 -16.280 ;
        RECT 26.760 -16.390 27.210 -16.280 ;
        RECT 24.910 -16.630 27.210 -16.390 ;
        RECT 24.910 -16.700 25.360 -16.630 ;
        RECT 8.160 -17.260 8.610 -17.210 ;
        RECT 6.520 -17.550 8.610 -17.260 ;
        RECT 6.520 -17.600 6.970 -17.550 ;
        RECT 1.420 -18.180 1.870 -18.080 ;
        RECT 2.260 -18.180 2.670 -17.750 ;
        RECT 5.420 -17.820 6.970 -17.600 ;
        RECT 7.350 -17.610 7.780 -17.550 ;
        RECT 8.160 -17.600 8.610 -17.550 ;
        RECT 9.210 -17.600 9.710 -17.210 ;
        RECT 8.160 -17.820 9.710 -17.600 ;
        RECT 18.920 -17.210 20.470 -16.990 ;
        RECT 18.920 -17.600 19.420 -17.210 ;
        RECT 20.020 -17.260 20.470 -17.210 ;
        RECT 20.850 -17.260 21.280 -17.200 ;
        RECT 21.660 -17.210 23.210 -16.990 ;
        RECT 25.960 -17.060 26.370 -16.630 ;
        RECT 26.760 -16.730 27.210 -16.630 ;
        RECT 28.420 -16.390 28.870 -16.280 ;
        RECT 30.270 -16.390 30.720 -16.280 ;
        RECT 28.420 -16.630 30.720 -16.390 ;
        RECT 28.420 -16.730 28.870 -16.630 ;
        RECT 29.260 -17.060 29.670 -16.630 ;
        RECT 30.270 -16.700 30.720 -16.630 ;
        RECT 31.670 -16.390 32.120 -16.310 ;
        RECT 32.720 -16.390 33.130 -15.950 ;
        RECT 33.520 -16.390 33.970 -16.280 ;
        RECT 31.670 -16.630 33.970 -16.390 ;
        RECT 31.670 -16.730 32.120 -16.630 ;
        RECT 33.520 -16.730 33.970 -16.630 ;
        RECT 35.160 -16.390 35.610 -16.280 ;
        RECT 36.000 -16.390 36.410 -15.950 ;
        RECT 39.180 -16.220 39.630 -15.940 ;
        RECT 43.000 -16.220 43.450 -15.940 ;
        RECT 52.680 -15.940 54.210 -15.730 ;
        RECT 54.590 -15.820 55.040 -15.730 ;
        RECT 55.420 -15.940 56.950 -15.730 ;
        RECT 37.010 -16.390 37.460 -16.310 ;
        RECT 35.160 -16.630 37.460 -16.390 ;
        RECT 35.160 -16.730 35.610 -16.630 ;
        RECT 37.010 -16.730 37.460 -16.630 ;
        RECT 38.410 -16.390 38.860 -16.280 ;
        RECT 40.260 -16.390 40.710 -16.280 ;
        RECT 38.410 -16.630 40.710 -16.390 ;
        RECT 38.410 -16.700 38.860 -16.630 ;
        RECT 21.660 -17.260 22.110 -17.210 ;
        RECT 20.020 -17.550 22.110 -17.260 ;
        RECT 20.020 -17.600 20.470 -17.550 ;
        RECT 3.270 -18.180 3.720 -18.110 ;
        RECT 1.420 -18.420 3.720 -18.180 ;
        RECT 1.420 -18.530 1.870 -18.420 ;
        RECT 3.270 -18.530 3.720 -18.420 ;
        RECT 4.670 -18.180 5.120 -18.080 ;
        RECT 6.520 -18.180 6.970 -18.080 ;
        RECT 4.670 -18.420 6.970 -18.180 ;
        RECT 4.670 -18.500 5.120 -18.420 ;
        RECT 5.720 -18.860 6.130 -18.420 ;
        RECT 6.520 -18.530 6.970 -18.420 ;
        RECT 8.160 -18.180 8.610 -18.080 ;
        RECT 10.010 -18.180 10.460 -18.080 ;
        RECT 8.160 -18.420 10.460 -18.180 ;
        RECT 8.160 -18.530 8.610 -18.420 ;
        RECT 9.000 -18.860 9.410 -18.420 ;
        RECT 10.010 -18.500 10.460 -18.420 ;
        RECT 11.410 -18.180 11.860 -18.110 ;
        RECT 12.460 -18.180 12.870 -17.750 ;
        RECT 13.260 -18.180 13.710 -18.080 ;
        RECT 11.410 -18.420 13.710 -18.180 ;
        RECT 11.410 -18.530 11.860 -18.420 ;
        RECT 13.260 -18.530 13.710 -18.420 ;
        RECT 14.920 -18.180 15.370 -18.080 ;
        RECT 15.760 -18.180 16.170 -17.750 ;
        RECT 18.920 -17.820 20.470 -17.600 ;
        RECT 20.850 -17.610 21.280 -17.550 ;
        RECT 21.660 -17.600 22.110 -17.550 ;
        RECT 22.710 -17.600 23.210 -17.210 ;
        RECT 21.660 -17.820 23.210 -17.600 ;
        RECT 32.420 -17.210 33.970 -16.990 ;
        RECT 32.420 -17.600 32.920 -17.210 ;
        RECT 33.520 -17.260 33.970 -17.210 ;
        RECT 34.350 -17.260 34.780 -17.200 ;
        RECT 35.160 -17.210 36.710 -16.990 ;
        RECT 39.460 -17.060 39.870 -16.630 ;
        RECT 40.260 -16.730 40.710 -16.630 ;
        RECT 41.920 -16.390 42.370 -16.280 ;
        RECT 43.770 -16.390 44.220 -16.280 ;
        RECT 41.920 -16.630 44.220 -16.390 ;
        RECT 41.920 -16.730 42.370 -16.630 ;
        RECT 42.760 -17.060 43.170 -16.630 ;
        RECT 43.770 -16.700 44.220 -16.630 ;
        RECT 45.170 -16.390 45.620 -16.310 ;
        RECT 46.220 -16.390 46.630 -15.950 ;
        RECT 47.020 -16.390 47.470 -16.280 ;
        RECT 45.170 -16.630 47.470 -16.390 ;
        RECT 45.170 -16.730 45.620 -16.630 ;
        RECT 47.020 -16.730 47.470 -16.630 ;
        RECT 48.660 -16.390 49.110 -16.280 ;
        RECT 49.500 -16.390 49.910 -15.950 ;
        RECT 52.680 -16.220 53.130 -15.940 ;
        RECT 56.500 -16.220 56.950 -15.940 ;
        RECT 66.180 -15.940 67.710 -15.730 ;
        RECT 68.090 -15.820 68.540 -15.730 ;
        RECT 68.920 -15.940 70.450 -15.730 ;
        RECT 50.510 -16.390 50.960 -16.310 ;
        RECT 48.660 -16.630 50.960 -16.390 ;
        RECT 48.660 -16.730 49.110 -16.630 ;
        RECT 50.510 -16.730 50.960 -16.630 ;
        RECT 51.910 -16.390 52.360 -16.280 ;
        RECT 53.760 -16.390 54.210 -16.280 ;
        RECT 51.910 -16.630 54.210 -16.390 ;
        RECT 51.910 -16.700 52.360 -16.630 ;
        RECT 35.160 -17.260 35.610 -17.210 ;
        RECT 33.520 -17.550 35.610 -17.260 ;
        RECT 33.520 -17.600 33.970 -17.550 ;
        RECT 16.770 -18.180 17.220 -18.110 ;
        RECT 14.920 -18.420 17.220 -18.180 ;
        RECT 14.920 -18.530 15.370 -18.420 ;
        RECT 16.770 -18.530 17.220 -18.420 ;
        RECT 18.170 -18.180 18.620 -18.080 ;
        RECT 20.020 -18.180 20.470 -18.080 ;
        RECT 18.170 -18.420 20.470 -18.180 ;
        RECT 18.170 -18.500 18.620 -18.420 ;
        RECT 12.180 -18.870 12.630 -18.590 ;
        RECT 16.000 -18.870 16.450 -18.590 ;
        RECT 19.220 -18.860 19.630 -18.420 ;
        RECT 20.020 -18.530 20.470 -18.420 ;
        RECT 21.660 -18.180 22.110 -18.080 ;
        RECT 23.510 -18.180 23.960 -18.080 ;
        RECT 21.660 -18.420 23.960 -18.180 ;
        RECT 21.660 -18.530 22.110 -18.420 ;
        RECT 22.500 -18.860 22.910 -18.420 ;
        RECT 23.510 -18.500 23.960 -18.420 ;
        RECT 24.910 -18.180 25.360 -18.110 ;
        RECT 25.960 -18.180 26.370 -17.750 ;
        RECT 26.760 -18.180 27.210 -18.080 ;
        RECT 24.910 -18.420 27.210 -18.180 ;
        RECT 24.910 -18.530 25.360 -18.420 ;
        RECT 26.760 -18.530 27.210 -18.420 ;
        RECT 28.420 -18.180 28.870 -18.080 ;
        RECT 29.260 -18.180 29.670 -17.750 ;
        RECT 32.420 -17.820 33.970 -17.600 ;
        RECT 34.350 -17.610 34.780 -17.550 ;
        RECT 35.160 -17.600 35.610 -17.550 ;
        RECT 36.210 -17.600 36.710 -17.210 ;
        RECT 35.160 -17.820 36.710 -17.600 ;
        RECT 45.920 -17.210 47.470 -16.990 ;
        RECT 45.920 -17.600 46.420 -17.210 ;
        RECT 47.020 -17.260 47.470 -17.210 ;
        RECT 47.850 -17.260 48.280 -17.200 ;
        RECT 48.660 -17.210 50.210 -16.990 ;
        RECT 52.960 -17.060 53.370 -16.630 ;
        RECT 53.760 -16.730 54.210 -16.630 ;
        RECT 55.420 -16.390 55.870 -16.280 ;
        RECT 57.270 -16.390 57.720 -16.280 ;
        RECT 55.420 -16.630 57.720 -16.390 ;
        RECT 55.420 -16.730 55.870 -16.630 ;
        RECT 56.260 -17.060 56.670 -16.630 ;
        RECT 57.270 -16.700 57.720 -16.630 ;
        RECT 58.670 -16.390 59.120 -16.310 ;
        RECT 59.720 -16.390 60.130 -15.950 ;
        RECT 60.520 -16.390 60.970 -16.280 ;
        RECT 58.670 -16.630 60.970 -16.390 ;
        RECT 58.670 -16.730 59.120 -16.630 ;
        RECT 60.520 -16.730 60.970 -16.630 ;
        RECT 62.160 -16.390 62.610 -16.280 ;
        RECT 63.000 -16.390 63.410 -15.950 ;
        RECT 66.180 -16.220 66.630 -15.940 ;
        RECT 70.000 -16.220 70.450 -15.940 ;
        RECT 79.680 -15.940 81.210 -15.730 ;
        RECT 81.590 -15.820 82.040 -15.730 ;
        RECT 82.420 -15.940 83.950 -15.730 ;
        RECT 64.010 -16.390 64.460 -16.310 ;
        RECT 62.160 -16.630 64.460 -16.390 ;
        RECT 62.160 -16.730 62.610 -16.630 ;
        RECT 64.010 -16.730 64.460 -16.630 ;
        RECT 65.410 -16.390 65.860 -16.280 ;
        RECT 67.260 -16.390 67.710 -16.280 ;
        RECT 65.410 -16.630 67.710 -16.390 ;
        RECT 65.410 -16.700 65.860 -16.630 ;
        RECT 48.660 -17.260 49.110 -17.210 ;
        RECT 47.020 -17.550 49.110 -17.260 ;
        RECT 47.020 -17.600 47.470 -17.550 ;
        RECT 30.270 -18.180 30.720 -18.110 ;
        RECT 28.420 -18.420 30.720 -18.180 ;
        RECT 28.420 -18.530 28.870 -18.420 ;
        RECT 30.270 -18.530 30.720 -18.420 ;
        RECT 31.670 -18.180 32.120 -18.080 ;
        RECT 33.520 -18.180 33.970 -18.080 ;
        RECT 31.670 -18.420 33.970 -18.180 ;
        RECT 31.670 -18.500 32.120 -18.420 ;
        RECT 12.180 -19.080 13.710 -18.870 ;
        RECT 14.090 -19.080 14.540 -18.990 ;
        RECT 14.920 -19.080 16.450 -18.870 ;
        RECT 25.680 -18.870 26.130 -18.590 ;
        RECT 29.500 -18.870 29.950 -18.590 ;
        RECT 32.720 -18.860 33.130 -18.420 ;
        RECT 33.520 -18.530 33.970 -18.420 ;
        RECT 35.160 -18.180 35.610 -18.080 ;
        RECT 37.010 -18.180 37.460 -18.080 ;
        RECT 35.160 -18.420 37.460 -18.180 ;
        RECT 35.160 -18.530 35.610 -18.420 ;
        RECT 36.000 -18.860 36.410 -18.420 ;
        RECT 37.010 -18.500 37.460 -18.420 ;
        RECT 38.410 -18.180 38.860 -18.110 ;
        RECT 39.460 -18.180 39.870 -17.750 ;
        RECT 40.260 -18.180 40.710 -18.080 ;
        RECT 38.410 -18.420 40.710 -18.180 ;
        RECT 38.410 -18.530 38.860 -18.420 ;
        RECT 40.260 -18.530 40.710 -18.420 ;
        RECT 41.920 -18.180 42.370 -18.080 ;
        RECT 42.760 -18.180 43.170 -17.750 ;
        RECT 45.920 -17.820 47.470 -17.600 ;
        RECT 47.850 -17.610 48.280 -17.550 ;
        RECT 48.660 -17.600 49.110 -17.550 ;
        RECT 49.710 -17.600 50.210 -17.210 ;
        RECT 48.660 -17.820 50.210 -17.600 ;
        RECT 59.420 -17.210 60.970 -16.990 ;
        RECT 59.420 -17.600 59.920 -17.210 ;
        RECT 60.520 -17.260 60.970 -17.210 ;
        RECT 61.350 -17.260 61.780 -17.200 ;
        RECT 62.160 -17.210 63.710 -16.990 ;
        RECT 66.460 -17.060 66.870 -16.630 ;
        RECT 67.260 -16.730 67.710 -16.630 ;
        RECT 68.920 -16.390 69.370 -16.280 ;
        RECT 70.770 -16.390 71.220 -16.280 ;
        RECT 68.920 -16.630 71.220 -16.390 ;
        RECT 68.920 -16.730 69.370 -16.630 ;
        RECT 69.760 -17.060 70.170 -16.630 ;
        RECT 70.770 -16.700 71.220 -16.630 ;
        RECT 72.170 -16.390 72.620 -16.310 ;
        RECT 73.220 -16.390 73.630 -15.950 ;
        RECT 74.020 -16.390 74.470 -16.280 ;
        RECT 72.170 -16.630 74.470 -16.390 ;
        RECT 72.170 -16.730 72.620 -16.630 ;
        RECT 74.020 -16.730 74.470 -16.630 ;
        RECT 75.660 -16.390 76.110 -16.280 ;
        RECT 76.500 -16.390 76.910 -15.950 ;
        RECT 79.680 -16.220 80.130 -15.940 ;
        RECT 83.500 -16.220 83.950 -15.940 ;
        RECT 93.180 -15.940 94.710 -15.730 ;
        RECT 95.090 -15.820 95.540 -15.730 ;
        RECT 95.920 -15.940 97.450 -15.730 ;
        RECT 77.510 -16.390 77.960 -16.310 ;
        RECT 75.660 -16.630 77.960 -16.390 ;
        RECT 75.660 -16.730 76.110 -16.630 ;
        RECT 77.510 -16.730 77.960 -16.630 ;
        RECT 78.910 -16.390 79.360 -16.280 ;
        RECT 80.760 -16.390 81.210 -16.280 ;
        RECT 78.910 -16.630 81.210 -16.390 ;
        RECT 78.910 -16.700 79.360 -16.630 ;
        RECT 62.160 -17.260 62.610 -17.210 ;
        RECT 60.520 -17.550 62.610 -17.260 ;
        RECT 60.520 -17.600 60.970 -17.550 ;
        RECT 43.770 -18.180 44.220 -18.110 ;
        RECT 41.920 -18.420 44.220 -18.180 ;
        RECT 41.920 -18.530 42.370 -18.420 ;
        RECT 43.770 -18.530 44.220 -18.420 ;
        RECT 45.170 -18.180 45.620 -18.080 ;
        RECT 47.020 -18.180 47.470 -18.080 ;
        RECT 45.170 -18.420 47.470 -18.180 ;
        RECT 45.170 -18.500 45.620 -18.420 ;
        RECT 25.680 -19.080 27.210 -18.870 ;
        RECT 27.590 -19.080 28.040 -18.990 ;
        RECT 28.420 -19.080 29.950 -18.870 ;
        RECT 39.180 -18.870 39.630 -18.590 ;
        RECT 43.000 -18.870 43.450 -18.590 ;
        RECT 46.220 -18.860 46.630 -18.420 ;
        RECT 47.020 -18.530 47.470 -18.420 ;
        RECT 48.660 -18.180 49.110 -18.080 ;
        RECT 50.510 -18.180 50.960 -18.080 ;
        RECT 48.660 -18.420 50.960 -18.180 ;
        RECT 48.660 -18.530 49.110 -18.420 ;
        RECT 49.500 -18.860 49.910 -18.420 ;
        RECT 50.510 -18.500 50.960 -18.420 ;
        RECT 51.910 -18.180 52.360 -18.110 ;
        RECT 52.960 -18.180 53.370 -17.750 ;
        RECT 53.760 -18.180 54.210 -18.080 ;
        RECT 51.910 -18.420 54.210 -18.180 ;
        RECT 51.910 -18.530 52.360 -18.420 ;
        RECT 53.760 -18.530 54.210 -18.420 ;
        RECT 55.420 -18.180 55.870 -18.080 ;
        RECT 56.260 -18.180 56.670 -17.750 ;
        RECT 59.420 -17.820 60.970 -17.600 ;
        RECT 61.350 -17.610 61.780 -17.550 ;
        RECT 62.160 -17.600 62.610 -17.550 ;
        RECT 63.210 -17.600 63.710 -17.210 ;
        RECT 62.160 -17.820 63.710 -17.600 ;
        RECT 72.920 -17.210 74.470 -16.990 ;
        RECT 72.920 -17.600 73.420 -17.210 ;
        RECT 74.020 -17.260 74.470 -17.210 ;
        RECT 74.850 -17.260 75.280 -17.200 ;
        RECT 75.660 -17.210 77.210 -16.990 ;
        RECT 79.960 -17.060 80.370 -16.630 ;
        RECT 80.760 -16.730 81.210 -16.630 ;
        RECT 82.420 -16.390 82.870 -16.280 ;
        RECT 84.270 -16.390 84.720 -16.280 ;
        RECT 82.420 -16.630 84.720 -16.390 ;
        RECT 82.420 -16.730 82.870 -16.630 ;
        RECT 83.260 -17.060 83.670 -16.630 ;
        RECT 84.270 -16.700 84.720 -16.630 ;
        RECT 85.670 -16.390 86.120 -16.310 ;
        RECT 86.720 -16.390 87.130 -15.950 ;
        RECT 87.520 -16.390 87.970 -16.280 ;
        RECT 85.670 -16.630 87.970 -16.390 ;
        RECT 85.670 -16.730 86.120 -16.630 ;
        RECT 87.520 -16.730 87.970 -16.630 ;
        RECT 89.160 -16.390 89.610 -16.280 ;
        RECT 90.000 -16.390 90.410 -15.950 ;
        RECT 93.180 -16.220 93.630 -15.940 ;
        RECT 97.000 -16.220 97.450 -15.940 ;
        RECT 106.680 -15.940 108.210 -15.730 ;
        RECT 108.590 -15.820 109.040 -15.730 ;
        RECT 109.420 -15.940 110.950 -15.730 ;
        RECT 91.010 -16.390 91.460 -16.310 ;
        RECT 89.160 -16.630 91.460 -16.390 ;
        RECT 89.160 -16.730 89.610 -16.630 ;
        RECT 91.010 -16.730 91.460 -16.630 ;
        RECT 92.410 -16.390 92.860 -16.280 ;
        RECT 94.260 -16.390 94.710 -16.280 ;
        RECT 92.410 -16.630 94.710 -16.390 ;
        RECT 92.410 -16.700 92.860 -16.630 ;
        RECT 75.660 -17.260 76.110 -17.210 ;
        RECT 74.020 -17.550 76.110 -17.260 ;
        RECT 74.020 -17.600 74.470 -17.550 ;
        RECT 57.270 -18.180 57.720 -18.110 ;
        RECT 55.420 -18.420 57.720 -18.180 ;
        RECT 55.420 -18.530 55.870 -18.420 ;
        RECT 57.270 -18.530 57.720 -18.420 ;
        RECT 58.670 -18.180 59.120 -18.080 ;
        RECT 60.520 -18.180 60.970 -18.080 ;
        RECT 58.670 -18.420 60.970 -18.180 ;
        RECT 58.670 -18.500 59.120 -18.420 ;
        RECT 39.180 -19.080 40.710 -18.870 ;
        RECT 41.090 -19.080 41.540 -18.990 ;
        RECT 41.920 -19.080 43.450 -18.870 ;
        RECT 52.680 -18.870 53.130 -18.590 ;
        RECT 56.500 -18.870 56.950 -18.590 ;
        RECT 59.720 -18.860 60.130 -18.420 ;
        RECT 60.520 -18.530 60.970 -18.420 ;
        RECT 62.160 -18.180 62.610 -18.080 ;
        RECT 64.010 -18.180 64.460 -18.080 ;
        RECT 62.160 -18.420 64.460 -18.180 ;
        RECT 62.160 -18.530 62.610 -18.420 ;
        RECT 63.000 -18.860 63.410 -18.420 ;
        RECT 64.010 -18.500 64.460 -18.420 ;
        RECT 65.410 -18.180 65.860 -18.110 ;
        RECT 66.460 -18.180 66.870 -17.750 ;
        RECT 67.260 -18.180 67.710 -18.080 ;
        RECT 65.410 -18.420 67.710 -18.180 ;
        RECT 65.410 -18.530 65.860 -18.420 ;
        RECT 67.260 -18.530 67.710 -18.420 ;
        RECT 68.920 -18.180 69.370 -18.080 ;
        RECT 69.760 -18.180 70.170 -17.750 ;
        RECT 72.920 -17.820 74.470 -17.600 ;
        RECT 74.850 -17.610 75.280 -17.550 ;
        RECT 75.660 -17.600 76.110 -17.550 ;
        RECT 76.710 -17.600 77.210 -17.210 ;
        RECT 75.660 -17.820 77.210 -17.600 ;
        RECT 86.420 -17.210 87.970 -16.990 ;
        RECT 86.420 -17.600 86.920 -17.210 ;
        RECT 87.520 -17.260 87.970 -17.210 ;
        RECT 88.350 -17.260 88.780 -17.200 ;
        RECT 89.160 -17.210 90.710 -16.990 ;
        RECT 93.460 -17.060 93.870 -16.630 ;
        RECT 94.260 -16.730 94.710 -16.630 ;
        RECT 95.920 -16.390 96.370 -16.280 ;
        RECT 97.770 -16.390 98.220 -16.280 ;
        RECT 95.920 -16.630 98.220 -16.390 ;
        RECT 95.920 -16.730 96.370 -16.630 ;
        RECT 96.760 -17.060 97.170 -16.630 ;
        RECT 97.770 -16.700 98.220 -16.630 ;
        RECT 99.170 -16.390 99.620 -16.310 ;
        RECT 100.220 -16.390 100.630 -15.950 ;
        RECT 101.020 -16.390 101.470 -16.280 ;
        RECT 99.170 -16.630 101.470 -16.390 ;
        RECT 99.170 -16.730 99.620 -16.630 ;
        RECT 101.020 -16.730 101.470 -16.630 ;
        RECT 102.660 -16.390 103.110 -16.280 ;
        RECT 103.500 -16.390 103.910 -15.950 ;
        RECT 106.680 -16.220 107.130 -15.940 ;
        RECT 110.500 -16.220 110.950 -15.940 ;
        RECT 120.180 -15.940 121.710 -15.730 ;
        RECT 122.090 -15.820 122.540 -15.730 ;
        RECT 122.920 -15.940 124.450 -15.730 ;
        RECT 104.510 -16.390 104.960 -16.310 ;
        RECT 102.660 -16.630 104.960 -16.390 ;
        RECT 102.660 -16.730 103.110 -16.630 ;
        RECT 104.510 -16.730 104.960 -16.630 ;
        RECT 105.910 -16.390 106.360 -16.280 ;
        RECT 107.760 -16.390 108.210 -16.280 ;
        RECT 105.910 -16.630 108.210 -16.390 ;
        RECT 105.910 -16.700 106.360 -16.630 ;
        RECT 89.160 -17.260 89.610 -17.210 ;
        RECT 87.520 -17.550 89.610 -17.260 ;
        RECT 87.520 -17.600 87.970 -17.550 ;
        RECT 70.770 -18.180 71.220 -18.110 ;
        RECT 68.920 -18.420 71.220 -18.180 ;
        RECT 68.920 -18.530 69.370 -18.420 ;
        RECT 70.770 -18.530 71.220 -18.420 ;
        RECT 72.170 -18.180 72.620 -18.080 ;
        RECT 74.020 -18.180 74.470 -18.080 ;
        RECT 72.170 -18.420 74.470 -18.180 ;
        RECT 72.170 -18.500 72.620 -18.420 ;
        RECT 52.680 -19.080 54.210 -18.870 ;
        RECT 54.590 -19.080 55.040 -18.990 ;
        RECT 55.420 -19.080 56.950 -18.870 ;
        RECT 66.180 -18.870 66.630 -18.590 ;
        RECT 70.000 -18.870 70.450 -18.590 ;
        RECT 73.220 -18.860 73.630 -18.420 ;
        RECT 74.020 -18.530 74.470 -18.420 ;
        RECT 75.660 -18.180 76.110 -18.080 ;
        RECT 77.510 -18.180 77.960 -18.080 ;
        RECT 75.660 -18.420 77.960 -18.180 ;
        RECT 75.660 -18.530 76.110 -18.420 ;
        RECT 76.500 -18.860 76.910 -18.420 ;
        RECT 77.510 -18.500 77.960 -18.420 ;
        RECT 78.910 -18.180 79.360 -18.110 ;
        RECT 79.960 -18.180 80.370 -17.750 ;
        RECT 80.760 -18.180 81.210 -18.080 ;
        RECT 78.910 -18.420 81.210 -18.180 ;
        RECT 78.910 -18.530 79.360 -18.420 ;
        RECT 80.760 -18.530 81.210 -18.420 ;
        RECT 82.420 -18.180 82.870 -18.080 ;
        RECT 83.260 -18.180 83.670 -17.750 ;
        RECT 86.420 -17.820 87.970 -17.600 ;
        RECT 88.350 -17.610 88.780 -17.550 ;
        RECT 89.160 -17.600 89.610 -17.550 ;
        RECT 90.210 -17.600 90.710 -17.210 ;
        RECT 89.160 -17.820 90.710 -17.600 ;
        RECT 99.920 -17.210 101.470 -16.990 ;
        RECT 99.920 -17.600 100.420 -17.210 ;
        RECT 101.020 -17.260 101.470 -17.210 ;
        RECT 101.850 -17.260 102.280 -17.200 ;
        RECT 102.660 -17.210 104.210 -16.990 ;
        RECT 106.960 -17.060 107.370 -16.630 ;
        RECT 107.760 -16.730 108.210 -16.630 ;
        RECT 109.420 -16.390 109.870 -16.280 ;
        RECT 111.270 -16.390 111.720 -16.280 ;
        RECT 109.420 -16.630 111.720 -16.390 ;
        RECT 109.420 -16.730 109.870 -16.630 ;
        RECT 110.260 -17.060 110.670 -16.630 ;
        RECT 111.270 -16.700 111.720 -16.630 ;
        RECT 112.670 -16.390 113.120 -16.310 ;
        RECT 113.720 -16.390 114.130 -15.950 ;
        RECT 114.520 -16.390 114.970 -16.280 ;
        RECT 112.670 -16.630 114.970 -16.390 ;
        RECT 112.670 -16.730 113.120 -16.630 ;
        RECT 114.520 -16.730 114.970 -16.630 ;
        RECT 116.160 -16.390 116.610 -16.280 ;
        RECT 117.000 -16.390 117.410 -15.950 ;
        RECT 120.180 -16.220 120.630 -15.940 ;
        RECT 124.000 -16.220 124.450 -15.940 ;
        RECT 133.680 -15.940 135.210 -15.730 ;
        RECT 135.590 -15.820 136.040 -15.730 ;
        RECT 136.420 -15.940 137.950 -15.730 ;
        RECT 118.010 -16.390 118.460 -16.310 ;
        RECT 116.160 -16.630 118.460 -16.390 ;
        RECT 116.160 -16.730 116.610 -16.630 ;
        RECT 118.010 -16.730 118.460 -16.630 ;
        RECT 119.410 -16.390 119.860 -16.280 ;
        RECT 121.260 -16.390 121.710 -16.280 ;
        RECT 119.410 -16.630 121.710 -16.390 ;
        RECT 119.410 -16.700 119.860 -16.630 ;
        RECT 102.660 -17.260 103.110 -17.210 ;
        RECT 101.020 -17.550 103.110 -17.260 ;
        RECT 101.020 -17.600 101.470 -17.550 ;
        RECT 84.270 -18.180 84.720 -18.110 ;
        RECT 82.420 -18.420 84.720 -18.180 ;
        RECT 82.420 -18.530 82.870 -18.420 ;
        RECT 84.270 -18.530 84.720 -18.420 ;
        RECT 85.670 -18.180 86.120 -18.080 ;
        RECT 87.520 -18.180 87.970 -18.080 ;
        RECT 85.670 -18.420 87.970 -18.180 ;
        RECT 85.670 -18.500 86.120 -18.420 ;
        RECT 66.180 -19.080 67.710 -18.870 ;
        RECT 68.090 -19.080 68.540 -18.990 ;
        RECT 68.920 -19.080 70.450 -18.870 ;
        RECT 79.680 -18.870 80.130 -18.590 ;
        RECT 83.500 -18.870 83.950 -18.590 ;
        RECT 86.720 -18.860 87.130 -18.420 ;
        RECT 87.520 -18.530 87.970 -18.420 ;
        RECT 89.160 -18.180 89.610 -18.080 ;
        RECT 91.010 -18.180 91.460 -18.080 ;
        RECT 89.160 -18.420 91.460 -18.180 ;
        RECT 89.160 -18.530 89.610 -18.420 ;
        RECT 90.000 -18.860 90.410 -18.420 ;
        RECT 91.010 -18.500 91.460 -18.420 ;
        RECT 92.410 -18.180 92.860 -18.110 ;
        RECT 93.460 -18.180 93.870 -17.750 ;
        RECT 94.260 -18.180 94.710 -18.080 ;
        RECT 92.410 -18.420 94.710 -18.180 ;
        RECT 92.410 -18.530 92.860 -18.420 ;
        RECT 94.260 -18.530 94.710 -18.420 ;
        RECT 95.920 -18.180 96.370 -18.080 ;
        RECT 96.760 -18.180 97.170 -17.750 ;
        RECT 99.920 -17.820 101.470 -17.600 ;
        RECT 101.850 -17.610 102.280 -17.550 ;
        RECT 102.660 -17.600 103.110 -17.550 ;
        RECT 103.710 -17.600 104.210 -17.210 ;
        RECT 102.660 -17.820 104.210 -17.600 ;
        RECT 113.420 -17.210 114.970 -16.990 ;
        RECT 113.420 -17.600 113.920 -17.210 ;
        RECT 114.520 -17.260 114.970 -17.210 ;
        RECT 115.350 -17.260 115.780 -17.200 ;
        RECT 116.160 -17.210 117.710 -16.990 ;
        RECT 120.460 -17.060 120.870 -16.630 ;
        RECT 121.260 -16.730 121.710 -16.630 ;
        RECT 122.920 -16.390 123.370 -16.280 ;
        RECT 124.770 -16.390 125.220 -16.280 ;
        RECT 122.920 -16.630 125.220 -16.390 ;
        RECT 122.920 -16.730 123.370 -16.630 ;
        RECT 123.760 -17.060 124.170 -16.630 ;
        RECT 124.770 -16.700 125.220 -16.630 ;
        RECT 126.170 -16.390 126.620 -16.310 ;
        RECT 127.220 -16.390 127.630 -15.950 ;
        RECT 128.020 -16.390 128.470 -16.280 ;
        RECT 126.170 -16.630 128.470 -16.390 ;
        RECT 126.170 -16.730 126.620 -16.630 ;
        RECT 128.020 -16.730 128.470 -16.630 ;
        RECT 129.660 -16.390 130.110 -16.280 ;
        RECT 130.500 -16.390 130.910 -15.950 ;
        RECT 133.680 -16.220 134.130 -15.940 ;
        RECT 137.500 -16.220 137.950 -15.940 ;
        RECT 147.180 -15.940 148.710 -15.730 ;
        RECT 149.090 -15.820 149.540 -15.730 ;
        RECT 149.920 -15.940 151.450 -15.730 ;
        RECT 131.510 -16.390 131.960 -16.310 ;
        RECT 129.660 -16.630 131.960 -16.390 ;
        RECT 129.660 -16.730 130.110 -16.630 ;
        RECT 131.510 -16.730 131.960 -16.630 ;
        RECT 132.910 -16.390 133.360 -16.280 ;
        RECT 134.760 -16.390 135.210 -16.280 ;
        RECT 132.910 -16.630 135.210 -16.390 ;
        RECT 132.910 -16.700 133.360 -16.630 ;
        RECT 116.160 -17.260 116.610 -17.210 ;
        RECT 114.520 -17.550 116.610 -17.260 ;
        RECT 114.520 -17.600 114.970 -17.550 ;
        RECT 97.770 -18.180 98.220 -18.110 ;
        RECT 95.920 -18.420 98.220 -18.180 ;
        RECT 95.920 -18.530 96.370 -18.420 ;
        RECT 97.770 -18.530 98.220 -18.420 ;
        RECT 99.170 -18.180 99.620 -18.080 ;
        RECT 101.020 -18.180 101.470 -18.080 ;
        RECT 99.170 -18.420 101.470 -18.180 ;
        RECT 99.170 -18.500 99.620 -18.420 ;
        RECT 79.680 -19.080 81.210 -18.870 ;
        RECT 81.590 -19.080 82.040 -18.990 ;
        RECT 82.420 -19.080 83.950 -18.870 ;
        RECT 93.180 -18.870 93.630 -18.590 ;
        RECT 97.000 -18.870 97.450 -18.590 ;
        RECT 100.220 -18.860 100.630 -18.420 ;
        RECT 101.020 -18.530 101.470 -18.420 ;
        RECT 102.660 -18.180 103.110 -18.080 ;
        RECT 104.510 -18.180 104.960 -18.080 ;
        RECT 102.660 -18.420 104.960 -18.180 ;
        RECT 102.660 -18.530 103.110 -18.420 ;
        RECT 103.500 -18.860 103.910 -18.420 ;
        RECT 104.510 -18.500 104.960 -18.420 ;
        RECT 105.910 -18.180 106.360 -18.110 ;
        RECT 106.960 -18.180 107.370 -17.750 ;
        RECT 107.760 -18.180 108.210 -18.080 ;
        RECT 105.910 -18.420 108.210 -18.180 ;
        RECT 105.910 -18.530 106.360 -18.420 ;
        RECT 107.760 -18.530 108.210 -18.420 ;
        RECT 109.420 -18.180 109.870 -18.080 ;
        RECT 110.260 -18.180 110.670 -17.750 ;
        RECT 113.420 -17.820 114.970 -17.600 ;
        RECT 115.350 -17.610 115.780 -17.550 ;
        RECT 116.160 -17.600 116.610 -17.550 ;
        RECT 117.210 -17.600 117.710 -17.210 ;
        RECT 116.160 -17.820 117.710 -17.600 ;
        RECT 126.920 -17.210 128.470 -16.990 ;
        RECT 126.920 -17.600 127.420 -17.210 ;
        RECT 128.020 -17.260 128.470 -17.210 ;
        RECT 128.850 -17.260 129.280 -17.200 ;
        RECT 129.660 -17.210 131.210 -16.990 ;
        RECT 133.960 -17.060 134.370 -16.630 ;
        RECT 134.760 -16.730 135.210 -16.630 ;
        RECT 136.420 -16.390 136.870 -16.280 ;
        RECT 138.270 -16.390 138.720 -16.280 ;
        RECT 136.420 -16.630 138.720 -16.390 ;
        RECT 136.420 -16.730 136.870 -16.630 ;
        RECT 137.260 -17.060 137.670 -16.630 ;
        RECT 138.270 -16.700 138.720 -16.630 ;
        RECT 139.670 -16.390 140.120 -16.310 ;
        RECT 140.720 -16.390 141.130 -15.950 ;
        RECT 141.520 -16.390 141.970 -16.280 ;
        RECT 139.670 -16.630 141.970 -16.390 ;
        RECT 139.670 -16.730 140.120 -16.630 ;
        RECT 141.520 -16.730 141.970 -16.630 ;
        RECT 143.160 -16.390 143.610 -16.280 ;
        RECT 144.000 -16.390 144.410 -15.950 ;
        RECT 147.180 -16.220 147.630 -15.940 ;
        RECT 151.000 -16.220 151.450 -15.940 ;
        RECT 160.680 -15.940 162.210 -15.730 ;
        RECT 162.590 -15.820 163.040 -15.730 ;
        RECT 163.420 -15.940 164.950 -15.730 ;
        RECT 145.010 -16.390 145.460 -16.310 ;
        RECT 143.160 -16.630 145.460 -16.390 ;
        RECT 143.160 -16.730 143.610 -16.630 ;
        RECT 145.010 -16.730 145.460 -16.630 ;
        RECT 146.410 -16.390 146.860 -16.280 ;
        RECT 148.260 -16.390 148.710 -16.280 ;
        RECT 146.410 -16.630 148.710 -16.390 ;
        RECT 146.410 -16.700 146.860 -16.630 ;
        RECT 129.660 -17.260 130.110 -17.210 ;
        RECT 128.020 -17.550 130.110 -17.260 ;
        RECT 128.020 -17.600 128.470 -17.550 ;
        RECT 111.270 -18.180 111.720 -18.110 ;
        RECT 109.420 -18.420 111.720 -18.180 ;
        RECT 109.420 -18.530 109.870 -18.420 ;
        RECT 111.270 -18.530 111.720 -18.420 ;
        RECT 112.670 -18.180 113.120 -18.080 ;
        RECT 114.520 -18.180 114.970 -18.080 ;
        RECT 112.670 -18.420 114.970 -18.180 ;
        RECT 112.670 -18.500 113.120 -18.420 ;
        RECT 93.180 -19.080 94.710 -18.870 ;
        RECT 95.090 -19.080 95.540 -18.990 ;
        RECT 95.920 -19.080 97.450 -18.870 ;
        RECT 106.680 -18.870 107.130 -18.590 ;
        RECT 110.500 -18.870 110.950 -18.590 ;
        RECT 113.720 -18.860 114.130 -18.420 ;
        RECT 114.520 -18.530 114.970 -18.420 ;
        RECT 116.160 -18.180 116.610 -18.080 ;
        RECT 118.010 -18.180 118.460 -18.080 ;
        RECT 116.160 -18.420 118.460 -18.180 ;
        RECT 116.160 -18.530 116.610 -18.420 ;
        RECT 117.000 -18.860 117.410 -18.420 ;
        RECT 118.010 -18.500 118.460 -18.420 ;
        RECT 119.410 -18.180 119.860 -18.110 ;
        RECT 120.460 -18.180 120.870 -17.750 ;
        RECT 121.260 -18.180 121.710 -18.080 ;
        RECT 119.410 -18.420 121.710 -18.180 ;
        RECT 119.410 -18.530 119.860 -18.420 ;
        RECT 121.260 -18.530 121.710 -18.420 ;
        RECT 122.920 -18.180 123.370 -18.080 ;
        RECT 123.760 -18.180 124.170 -17.750 ;
        RECT 126.920 -17.820 128.470 -17.600 ;
        RECT 128.850 -17.610 129.280 -17.550 ;
        RECT 129.660 -17.600 130.110 -17.550 ;
        RECT 130.710 -17.600 131.210 -17.210 ;
        RECT 129.660 -17.820 131.210 -17.600 ;
        RECT 140.420 -17.210 141.970 -16.990 ;
        RECT 140.420 -17.600 140.920 -17.210 ;
        RECT 141.520 -17.260 141.970 -17.210 ;
        RECT 142.350 -17.260 142.780 -17.200 ;
        RECT 143.160 -17.210 144.710 -16.990 ;
        RECT 147.460 -17.060 147.870 -16.630 ;
        RECT 148.260 -16.730 148.710 -16.630 ;
        RECT 149.920 -16.390 150.370 -16.280 ;
        RECT 151.770 -16.390 152.220 -16.280 ;
        RECT 149.920 -16.630 152.220 -16.390 ;
        RECT 149.920 -16.730 150.370 -16.630 ;
        RECT 150.760 -17.060 151.170 -16.630 ;
        RECT 151.770 -16.700 152.220 -16.630 ;
        RECT 153.170 -16.390 153.620 -16.310 ;
        RECT 154.220 -16.390 154.630 -15.950 ;
        RECT 155.020 -16.390 155.470 -16.280 ;
        RECT 153.170 -16.630 155.470 -16.390 ;
        RECT 153.170 -16.730 153.620 -16.630 ;
        RECT 155.020 -16.730 155.470 -16.630 ;
        RECT 156.660 -16.390 157.110 -16.280 ;
        RECT 157.500 -16.390 157.910 -15.950 ;
        RECT 160.680 -16.220 161.130 -15.940 ;
        RECT 164.500 -16.220 164.950 -15.940 ;
        RECT 174.180 -15.940 175.710 -15.730 ;
        RECT 176.090 -15.820 176.540 -15.730 ;
        RECT 176.920 -15.940 178.450 -15.730 ;
        RECT 158.510 -16.390 158.960 -16.310 ;
        RECT 156.660 -16.630 158.960 -16.390 ;
        RECT 156.660 -16.730 157.110 -16.630 ;
        RECT 158.510 -16.730 158.960 -16.630 ;
        RECT 159.910 -16.390 160.360 -16.280 ;
        RECT 161.760 -16.390 162.210 -16.280 ;
        RECT 159.910 -16.630 162.210 -16.390 ;
        RECT 159.910 -16.700 160.360 -16.630 ;
        RECT 143.160 -17.260 143.610 -17.210 ;
        RECT 141.520 -17.550 143.610 -17.260 ;
        RECT 141.520 -17.600 141.970 -17.550 ;
        RECT 124.770 -18.180 125.220 -18.110 ;
        RECT 122.920 -18.420 125.220 -18.180 ;
        RECT 122.920 -18.530 123.370 -18.420 ;
        RECT 124.770 -18.530 125.220 -18.420 ;
        RECT 126.170 -18.180 126.620 -18.080 ;
        RECT 128.020 -18.180 128.470 -18.080 ;
        RECT 126.170 -18.420 128.470 -18.180 ;
        RECT 126.170 -18.500 126.620 -18.420 ;
        RECT 106.680 -19.080 108.210 -18.870 ;
        RECT 108.590 -19.080 109.040 -18.990 ;
        RECT 109.420 -19.080 110.950 -18.870 ;
        RECT 120.180 -18.870 120.630 -18.590 ;
        RECT 124.000 -18.870 124.450 -18.590 ;
        RECT 127.220 -18.860 127.630 -18.420 ;
        RECT 128.020 -18.530 128.470 -18.420 ;
        RECT 129.660 -18.180 130.110 -18.080 ;
        RECT 131.510 -18.180 131.960 -18.080 ;
        RECT 129.660 -18.420 131.960 -18.180 ;
        RECT 129.660 -18.530 130.110 -18.420 ;
        RECT 130.500 -18.860 130.910 -18.420 ;
        RECT 131.510 -18.500 131.960 -18.420 ;
        RECT 132.910 -18.180 133.360 -18.110 ;
        RECT 133.960 -18.180 134.370 -17.750 ;
        RECT 134.760 -18.180 135.210 -18.080 ;
        RECT 132.910 -18.420 135.210 -18.180 ;
        RECT 132.910 -18.530 133.360 -18.420 ;
        RECT 134.760 -18.530 135.210 -18.420 ;
        RECT 136.420 -18.180 136.870 -18.080 ;
        RECT 137.260 -18.180 137.670 -17.750 ;
        RECT 140.420 -17.820 141.970 -17.600 ;
        RECT 142.350 -17.610 142.780 -17.550 ;
        RECT 143.160 -17.600 143.610 -17.550 ;
        RECT 144.210 -17.600 144.710 -17.210 ;
        RECT 143.160 -17.820 144.710 -17.600 ;
        RECT 153.920 -17.210 155.470 -16.990 ;
        RECT 153.920 -17.600 154.420 -17.210 ;
        RECT 155.020 -17.260 155.470 -17.210 ;
        RECT 155.850 -17.260 156.280 -17.200 ;
        RECT 156.660 -17.210 158.210 -16.990 ;
        RECT 160.960 -17.060 161.370 -16.630 ;
        RECT 161.760 -16.730 162.210 -16.630 ;
        RECT 163.420 -16.390 163.870 -16.280 ;
        RECT 165.270 -16.390 165.720 -16.280 ;
        RECT 163.420 -16.630 165.720 -16.390 ;
        RECT 163.420 -16.730 163.870 -16.630 ;
        RECT 164.260 -17.060 164.670 -16.630 ;
        RECT 165.270 -16.700 165.720 -16.630 ;
        RECT 166.670 -16.390 167.120 -16.310 ;
        RECT 167.720 -16.390 168.130 -15.950 ;
        RECT 168.520 -16.390 168.970 -16.280 ;
        RECT 166.670 -16.630 168.970 -16.390 ;
        RECT 166.670 -16.730 167.120 -16.630 ;
        RECT 168.520 -16.730 168.970 -16.630 ;
        RECT 170.160 -16.390 170.610 -16.280 ;
        RECT 171.000 -16.390 171.410 -15.950 ;
        RECT 174.180 -16.220 174.630 -15.940 ;
        RECT 178.000 -16.220 178.450 -15.940 ;
        RECT 187.680 -15.940 189.210 -15.730 ;
        RECT 189.590 -15.820 190.040 -15.730 ;
        RECT 190.420 -15.940 191.950 -15.730 ;
        RECT 172.010 -16.390 172.460 -16.310 ;
        RECT 170.160 -16.630 172.460 -16.390 ;
        RECT 170.160 -16.730 170.610 -16.630 ;
        RECT 172.010 -16.730 172.460 -16.630 ;
        RECT 173.410 -16.390 173.860 -16.280 ;
        RECT 175.260 -16.390 175.710 -16.280 ;
        RECT 173.410 -16.630 175.710 -16.390 ;
        RECT 173.410 -16.700 173.860 -16.630 ;
        RECT 156.660 -17.260 157.110 -17.210 ;
        RECT 155.020 -17.550 157.110 -17.260 ;
        RECT 155.020 -17.600 155.470 -17.550 ;
        RECT 138.270 -18.180 138.720 -18.110 ;
        RECT 136.420 -18.420 138.720 -18.180 ;
        RECT 136.420 -18.530 136.870 -18.420 ;
        RECT 138.270 -18.530 138.720 -18.420 ;
        RECT 139.670 -18.180 140.120 -18.080 ;
        RECT 141.520 -18.180 141.970 -18.080 ;
        RECT 139.670 -18.420 141.970 -18.180 ;
        RECT 139.670 -18.500 140.120 -18.420 ;
        RECT 120.180 -19.080 121.710 -18.870 ;
        RECT 122.090 -19.080 122.540 -18.990 ;
        RECT 122.920 -19.080 124.450 -18.870 ;
        RECT 133.680 -18.870 134.130 -18.590 ;
        RECT 137.500 -18.870 137.950 -18.590 ;
        RECT 140.720 -18.860 141.130 -18.420 ;
        RECT 141.520 -18.530 141.970 -18.420 ;
        RECT 143.160 -18.180 143.610 -18.080 ;
        RECT 145.010 -18.180 145.460 -18.080 ;
        RECT 143.160 -18.420 145.460 -18.180 ;
        RECT 143.160 -18.530 143.610 -18.420 ;
        RECT 144.000 -18.860 144.410 -18.420 ;
        RECT 145.010 -18.500 145.460 -18.420 ;
        RECT 146.410 -18.180 146.860 -18.110 ;
        RECT 147.460 -18.180 147.870 -17.750 ;
        RECT 148.260 -18.180 148.710 -18.080 ;
        RECT 146.410 -18.420 148.710 -18.180 ;
        RECT 146.410 -18.530 146.860 -18.420 ;
        RECT 148.260 -18.530 148.710 -18.420 ;
        RECT 149.920 -18.180 150.370 -18.080 ;
        RECT 150.760 -18.180 151.170 -17.750 ;
        RECT 153.920 -17.820 155.470 -17.600 ;
        RECT 155.850 -17.610 156.280 -17.550 ;
        RECT 156.660 -17.600 157.110 -17.550 ;
        RECT 157.710 -17.600 158.210 -17.210 ;
        RECT 156.660 -17.820 158.210 -17.600 ;
        RECT 167.420 -17.210 168.970 -16.990 ;
        RECT 167.420 -17.600 167.920 -17.210 ;
        RECT 168.520 -17.260 168.970 -17.210 ;
        RECT 169.350 -17.260 169.780 -17.200 ;
        RECT 170.160 -17.210 171.710 -16.990 ;
        RECT 174.460 -17.060 174.870 -16.630 ;
        RECT 175.260 -16.730 175.710 -16.630 ;
        RECT 176.920 -16.390 177.370 -16.280 ;
        RECT 178.770 -16.390 179.220 -16.280 ;
        RECT 176.920 -16.630 179.220 -16.390 ;
        RECT 176.920 -16.730 177.370 -16.630 ;
        RECT 177.760 -17.060 178.170 -16.630 ;
        RECT 178.770 -16.700 179.220 -16.630 ;
        RECT 180.170 -16.390 180.620 -16.310 ;
        RECT 181.220 -16.390 181.630 -15.950 ;
        RECT 182.020 -16.390 182.470 -16.280 ;
        RECT 180.170 -16.630 182.470 -16.390 ;
        RECT 180.170 -16.730 180.620 -16.630 ;
        RECT 182.020 -16.730 182.470 -16.630 ;
        RECT 183.660 -16.390 184.110 -16.280 ;
        RECT 184.500 -16.390 184.910 -15.950 ;
        RECT 187.680 -16.220 188.130 -15.940 ;
        RECT 191.500 -16.220 191.950 -15.940 ;
        RECT 201.180 -15.940 202.710 -15.730 ;
        RECT 203.090 -15.820 203.540 -15.730 ;
        RECT 203.920 -15.940 205.450 -15.730 ;
        RECT 185.510 -16.390 185.960 -16.310 ;
        RECT 183.660 -16.630 185.960 -16.390 ;
        RECT 183.660 -16.730 184.110 -16.630 ;
        RECT 185.510 -16.730 185.960 -16.630 ;
        RECT 186.910 -16.390 187.360 -16.280 ;
        RECT 188.760 -16.390 189.210 -16.280 ;
        RECT 186.910 -16.630 189.210 -16.390 ;
        RECT 186.910 -16.700 187.360 -16.630 ;
        RECT 170.160 -17.260 170.610 -17.210 ;
        RECT 168.520 -17.550 170.610 -17.260 ;
        RECT 168.520 -17.600 168.970 -17.550 ;
        RECT 151.770 -18.180 152.220 -18.110 ;
        RECT 149.920 -18.420 152.220 -18.180 ;
        RECT 149.920 -18.530 150.370 -18.420 ;
        RECT 151.770 -18.530 152.220 -18.420 ;
        RECT 153.170 -18.180 153.620 -18.080 ;
        RECT 155.020 -18.180 155.470 -18.080 ;
        RECT 153.170 -18.420 155.470 -18.180 ;
        RECT 153.170 -18.500 153.620 -18.420 ;
        RECT 133.680 -19.080 135.210 -18.870 ;
        RECT 135.590 -19.080 136.040 -18.990 ;
        RECT 136.420 -19.080 137.950 -18.870 ;
        RECT 147.180 -18.870 147.630 -18.590 ;
        RECT 151.000 -18.870 151.450 -18.590 ;
        RECT 154.220 -18.860 154.630 -18.420 ;
        RECT 155.020 -18.530 155.470 -18.420 ;
        RECT 156.660 -18.180 157.110 -18.080 ;
        RECT 158.510 -18.180 158.960 -18.080 ;
        RECT 156.660 -18.420 158.960 -18.180 ;
        RECT 156.660 -18.530 157.110 -18.420 ;
        RECT 157.500 -18.860 157.910 -18.420 ;
        RECT 158.510 -18.500 158.960 -18.420 ;
        RECT 159.910 -18.180 160.360 -18.110 ;
        RECT 160.960 -18.180 161.370 -17.750 ;
        RECT 161.760 -18.180 162.210 -18.080 ;
        RECT 159.910 -18.420 162.210 -18.180 ;
        RECT 159.910 -18.530 160.360 -18.420 ;
        RECT 161.760 -18.530 162.210 -18.420 ;
        RECT 163.420 -18.180 163.870 -18.080 ;
        RECT 164.260 -18.180 164.670 -17.750 ;
        RECT 167.420 -17.820 168.970 -17.600 ;
        RECT 169.350 -17.610 169.780 -17.550 ;
        RECT 170.160 -17.600 170.610 -17.550 ;
        RECT 171.210 -17.600 171.710 -17.210 ;
        RECT 170.160 -17.820 171.710 -17.600 ;
        RECT 180.920 -17.210 182.470 -16.990 ;
        RECT 180.920 -17.600 181.420 -17.210 ;
        RECT 182.020 -17.260 182.470 -17.210 ;
        RECT 182.850 -17.260 183.280 -17.200 ;
        RECT 183.660 -17.210 185.210 -16.990 ;
        RECT 187.960 -17.060 188.370 -16.630 ;
        RECT 188.760 -16.730 189.210 -16.630 ;
        RECT 190.420 -16.390 190.870 -16.280 ;
        RECT 192.270 -16.390 192.720 -16.280 ;
        RECT 190.420 -16.630 192.720 -16.390 ;
        RECT 190.420 -16.730 190.870 -16.630 ;
        RECT 191.260 -17.060 191.670 -16.630 ;
        RECT 192.270 -16.700 192.720 -16.630 ;
        RECT 193.670 -16.390 194.120 -16.310 ;
        RECT 194.720 -16.390 195.130 -15.950 ;
        RECT 195.520 -16.390 195.970 -16.280 ;
        RECT 193.670 -16.630 195.970 -16.390 ;
        RECT 193.670 -16.730 194.120 -16.630 ;
        RECT 195.520 -16.730 195.970 -16.630 ;
        RECT 197.160 -16.390 197.610 -16.280 ;
        RECT 198.000 -16.390 198.410 -15.950 ;
        RECT 201.180 -16.220 201.630 -15.940 ;
        RECT 205.000 -16.220 205.450 -15.940 ;
        RECT 214.680 -15.940 216.210 -15.730 ;
        RECT 216.590 -15.820 217.030 -15.730 ;
        RECT 199.010 -16.390 199.460 -16.310 ;
        RECT 197.160 -16.630 199.460 -16.390 ;
        RECT 197.160 -16.730 197.610 -16.630 ;
        RECT 199.010 -16.730 199.460 -16.630 ;
        RECT 200.410 -16.390 200.860 -16.280 ;
        RECT 202.260 -16.390 202.710 -16.280 ;
        RECT 200.410 -16.630 202.710 -16.390 ;
        RECT 200.410 -16.700 200.860 -16.630 ;
        RECT 183.660 -17.260 184.110 -17.210 ;
        RECT 182.020 -17.550 184.110 -17.260 ;
        RECT 182.020 -17.600 182.470 -17.550 ;
        RECT 165.270 -18.180 165.720 -18.110 ;
        RECT 163.420 -18.420 165.720 -18.180 ;
        RECT 163.420 -18.530 163.870 -18.420 ;
        RECT 165.270 -18.530 165.720 -18.420 ;
        RECT 166.670 -18.180 167.120 -18.080 ;
        RECT 168.520 -18.180 168.970 -18.080 ;
        RECT 166.670 -18.420 168.970 -18.180 ;
        RECT 166.670 -18.500 167.120 -18.420 ;
        RECT 147.180 -19.080 148.710 -18.870 ;
        RECT 149.090 -19.080 149.540 -18.990 ;
        RECT 149.920 -19.080 151.450 -18.870 ;
        RECT 160.680 -18.870 161.130 -18.590 ;
        RECT 164.500 -18.870 164.950 -18.590 ;
        RECT 167.720 -18.860 168.130 -18.420 ;
        RECT 168.520 -18.530 168.970 -18.420 ;
        RECT 170.160 -18.180 170.610 -18.080 ;
        RECT 172.010 -18.180 172.460 -18.080 ;
        RECT 170.160 -18.420 172.460 -18.180 ;
        RECT 170.160 -18.530 170.610 -18.420 ;
        RECT 171.000 -18.860 171.410 -18.420 ;
        RECT 172.010 -18.500 172.460 -18.420 ;
        RECT 173.410 -18.180 173.860 -18.110 ;
        RECT 174.460 -18.180 174.870 -17.750 ;
        RECT 175.260 -18.180 175.710 -18.080 ;
        RECT 173.410 -18.420 175.710 -18.180 ;
        RECT 173.410 -18.530 173.860 -18.420 ;
        RECT 175.260 -18.530 175.710 -18.420 ;
        RECT 176.920 -18.180 177.370 -18.080 ;
        RECT 177.760 -18.180 178.170 -17.750 ;
        RECT 180.920 -17.820 182.470 -17.600 ;
        RECT 182.850 -17.610 183.280 -17.550 ;
        RECT 183.660 -17.600 184.110 -17.550 ;
        RECT 184.710 -17.600 185.210 -17.210 ;
        RECT 183.660 -17.820 185.210 -17.600 ;
        RECT 194.420 -17.210 195.970 -16.990 ;
        RECT 194.420 -17.600 194.920 -17.210 ;
        RECT 195.520 -17.260 195.970 -17.210 ;
        RECT 196.350 -17.260 196.780 -17.200 ;
        RECT 197.160 -17.210 198.710 -16.990 ;
        RECT 201.460 -17.060 201.870 -16.630 ;
        RECT 202.260 -16.730 202.710 -16.630 ;
        RECT 203.920 -16.390 204.370 -16.280 ;
        RECT 205.770 -16.390 206.220 -16.280 ;
        RECT 203.920 -16.630 206.220 -16.390 ;
        RECT 203.920 -16.730 204.370 -16.630 ;
        RECT 204.760 -17.060 205.170 -16.630 ;
        RECT 205.770 -16.700 206.220 -16.630 ;
        RECT 207.170 -16.390 207.620 -16.310 ;
        RECT 208.220 -16.390 208.630 -15.950 ;
        RECT 209.020 -16.390 209.470 -16.280 ;
        RECT 207.170 -16.630 209.470 -16.390 ;
        RECT 207.170 -16.730 207.620 -16.630 ;
        RECT 209.020 -16.730 209.470 -16.630 ;
        RECT 210.660 -16.390 211.110 -16.280 ;
        RECT 211.500 -16.390 211.910 -15.950 ;
        RECT 214.680 -16.220 215.130 -15.940 ;
        RECT 212.510 -16.390 212.960 -16.310 ;
        RECT 210.660 -16.630 212.960 -16.390 ;
        RECT 210.660 -16.730 211.110 -16.630 ;
        RECT 212.510 -16.730 212.960 -16.630 ;
        RECT 213.910 -16.390 214.360 -16.280 ;
        RECT 215.760 -16.390 216.210 -16.280 ;
        RECT 213.910 -16.630 216.210 -16.390 ;
        RECT 213.910 -16.700 214.360 -16.630 ;
        RECT 197.160 -17.260 197.610 -17.210 ;
        RECT 195.520 -17.550 197.610 -17.260 ;
        RECT 195.520 -17.600 195.970 -17.550 ;
        RECT 178.770 -18.180 179.220 -18.110 ;
        RECT 176.920 -18.420 179.220 -18.180 ;
        RECT 176.920 -18.530 177.370 -18.420 ;
        RECT 178.770 -18.530 179.220 -18.420 ;
        RECT 180.170 -18.180 180.620 -18.080 ;
        RECT 182.020 -18.180 182.470 -18.080 ;
        RECT 180.170 -18.420 182.470 -18.180 ;
        RECT 180.170 -18.500 180.620 -18.420 ;
        RECT 160.680 -19.080 162.210 -18.870 ;
        RECT 162.590 -19.080 163.040 -18.990 ;
        RECT 163.420 -19.080 164.950 -18.870 ;
        RECT 174.180 -18.870 174.630 -18.590 ;
        RECT 178.000 -18.870 178.450 -18.590 ;
        RECT 181.220 -18.860 181.630 -18.420 ;
        RECT 182.020 -18.530 182.470 -18.420 ;
        RECT 183.660 -18.180 184.110 -18.080 ;
        RECT 185.510 -18.180 185.960 -18.080 ;
        RECT 183.660 -18.420 185.960 -18.180 ;
        RECT 183.660 -18.530 184.110 -18.420 ;
        RECT 184.500 -18.860 184.910 -18.420 ;
        RECT 185.510 -18.500 185.960 -18.420 ;
        RECT 186.910 -18.180 187.360 -18.110 ;
        RECT 187.960 -18.180 188.370 -17.750 ;
        RECT 188.760 -18.180 189.210 -18.080 ;
        RECT 186.910 -18.420 189.210 -18.180 ;
        RECT 186.910 -18.530 187.360 -18.420 ;
        RECT 188.760 -18.530 189.210 -18.420 ;
        RECT 190.420 -18.180 190.870 -18.080 ;
        RECT 191.260 -18.180 191.670 -17.750 ;
        RECT 194.420 -17.820 195.970 -17.600 ;
        RECT 196.350 -17.610 196.780 -17.550 ;
        RECT 197.160 -17.600 197.610 -17.550 ;
        RECT 198.210 -17.600 198.710 -17.210 ;
        RECT 197.160 -17.820 198.710 -17.600 ;
        RECT 207.920 -17.210 209.470 -16.990 ;
        RECT 207.920 -17.600 208.420 -17.210 ;
        RECT 209.020 -17.260 209.470 -17.210 ;
        RECT 209.850 -17.260 210.280 -17.200 ;
        RECT 210.660 -17.210 212.210 -16.990 ;
        RECT 214.960 -17.060 215.370 -16.630 ;
        RECT 215.760 -16.730 216.210 -16.630 ;
        RECT 210.660 -17.260 211.110 -17.210 ;
        RECT 209.020 -17.550 211.110 -17.260 ;
        RECT 209.020 -17.600 209.470 -17.550 ;
        RECT 192.270 -18.180 192.720 -18.110 ;
        RECT 190.420 -18.420 192.720 -18.180 ;
        RECT 190.420 -18.530 190.870 -18.420 ;
        RECT 192.270 -18.530 192.720 -18.420 ;
        RECT 193.670 -18.180 194.120 -18.080 ;
        RECT 195.520 -18.180 195.970 -18.080 ;
        RECT 193.670 -18.420 195.970 -18.180 ;
        RECT 193.670 -18.500 194.120 -18.420 ;
        RECT 174.180 -19.080 175.710 -18.870 ;
        RECT 176.090 -19.080 176.540 -18.990 ;
        RECT 176.920 -19.080 178.450 -18.870 ;
        RECT 187.680 -18.870 188.130 -18.590 ;
        RECT 191.500 -18.870 191.950 -18.590 ;
        RECT 194.720 -18.860 195.130 -18.420 ;
        RECT 195.520 -18.530 195.970 -18.420 ;
        RECT 197.160 -18.180 197.610 -18.080 ;
        RECT 199.010 -18.180 199.460 -18.080 ;
        RECT 197.160 -18.420 199.460 -18.180 ;
        RECT 197.160 -18.530 197.610 -18.420 ;
        RECT 198.000 -18.860 198.410 -18.420 ;
        RECT 199.010 -18.500 199.460 -18.420 ;
        RECT 200.410 -18.180 200.860 -18.110 ;
        RECT 201.460 -18.180 201.870 -17.750 ;
        RECT 202.260 -18.180 202.710 -18.080 ;
        RECT 200.410 -18.420 202.710 -18.180 ;
        RECT 200.410 -18.530 200.860 -18.420 ;
        RECT 202.260 -18.530 202.710 -18.420 ;
        RECT 203.920 -18.180 204.370 -18.080 ;
        RECT 204.760 -18.180 205.170 -17.750 ;
        RECT 207.920 -17.820 209.470 -17.600 ;
        RECT 209.850 -17.610 210.280 -17.550 ;
        RECT 210.660 -17.600 211.110 -17.550 ;
        RECT 211.710 -17.600 212.210 -17.210 ;
        RECT 210.660 -17.820 212.210 -17.600 ;
        RECT 205.770 -18.180 206.220 -18.110 ;
        RECT 203.920 -18.420 206.220 -18.180 ;
        RECT 203.920 -18.530 204.370 -18.420 ;
        RECT 205.770 -18.530 206.220 -18.420 ;
        RECT 207.170 -18.180 207.620 -18.080 ;
        RECT 209.020 -18.180 209.470 -18.080 ;
        RECT 207.170 -18.420 209.470 -18.180 ;
        RECT 207.170 -18.500 207.620 -18.420 ;
        RECT 187.680 -19.080 189.210 -18.870 ;
        RECT 189.590 -19.080 190.040 -18.990 ;
        RECT 190.420 -19.080 191.950 -18.870 ;
        RECT 201.180 -18.870 201.630 -18.590 ;
        RECT 205.000 -18.870 205.450 -18.590 ;
        RECT 208.220 -18.860 208.630 -18.420 ;
        RECT 209.020 -18.530 209.470 -18.420 ;
        RECT 210.660 -18.180 211.110 -18.080 ;
        RECT 212.510 -18.180 212.960 -18.080 ;
        RECT 210.660 -18.420 212.960 -18.180 ;
        RECT 210.660 -18.530 211.110 -18.420 ;
        RECT 211.500 -18.860 211.910 -18.420 ;
        RECT 212.510 -18.500 212.960 -18.420 ;
        RECT 213.910 -18.180 214.360 -18.110 ;
        RECT 214.960 -18.180 215.370 -17.750 ;
        RECT 215.760 -18.180 216.210 -18.080 ;
        RECT 213.910 -18.420 216.210 -18.180 ;
        RECT 213.910 -18.530 214.360 -18.420 ;
        RECT 215.760 -18.530 216.210 -18.420 ;
        RECT 201.180 -19.080 202.710 -18.870 ;
        RECT 203.090 -19.080 203.540 -18.990 ;
        RECT 203.920 -19.080 205.450 -18.870 ;
        RECT 214.680 -18.870 215.130 -18.590 ;
        RECT 214.680 -19.080 216.210 -18.870 ;
        RECT 216.590 -19.080 217.030 -18.990 ;
        RECT 13.260 -19.340 15.370 -19.080 ;
        RECT 26.760 -19.340 28.870 -19.080 ;
        RECT 40.260 -19.340 42.370 -19.080 ;
        RECT 53.760 -19.340 55.870 -19.080 ;
        RECT 67.260 -19.340 69.370 -19.080 ;
        RECT 80.760 -19.340 82.870 -19.080 ;
        RECT 94.260 -19.340 96.370 -19.080 ;
        RECT 107.760 -19.340 109.870 -19.080 ;
        RECT 121.260 -19.340 123.370 -19.080 ;
        RECT 134.760 -19.340 136.870 -19.080 ;
        RECT 148.260 -19.340 150.370 -19.080 ;
        RECT 161.760 -19.340 163.870 -19.080 ;
        RECT 175.260 -19.340 177.370 -19.080 ;
        RECT 188.760 -19.340 190.870 -19.080 ;
        RECT 202.260 -19.340 204.370 -19.080 ;
        RECT 215.760 -19.340 217.030 -19.080 ;
        RECT 12.180 -19.550 13.710 -19.340 ;
        RECT 14.090 -19.430 14.540 -19.340 ;
        RECT 14.920 -19.550 16.450 -19.340 ;
        RECT 1.420 -20.000 1.870 -19.890 ;
        RECT 3.270 -20.000 3.720 -19.890 ;
        RECT 1.420 -20.240 3.720 -20.000 ;
        RECT 1.420 -20.340 1.870 -20.240 ;
        RECT 2.260 -20.670 2.670 -20.240 ;
        RECT 3.270 -20.310 3.720 -20.240 ;
        RECT 4.670 -20.000 5.120 -19.920 ;
        RECT 5.720 -20.000 6.130 -19.560 ;
        RECT 6.520 -20.000 6.970 -19.890 ;
        RECT 4.670 -20.240 6.970 -20.000 ;
        RECT 4.670 -20.340 5.120 -20.240 ;
        RECT 6.520 -20.340 6.970 -20.240 ;
        RECT 8.160 -20.000 8.610 -19.890 ;
        RECT 9.000 -20.000 9.410 -19.560 ;
        RECT 12.180 -19.830 12.630 -19.550 ;
        RECT 16.000 -19.830 16.450 -19.550 ;
        RECT 25.680 -19.550 27.210 -19.340 ;
        RECT 27.590 -19.430 28.040 -19.340 ;
        RECT 28.420 -19.550 29.950 -19.340 ;
        RECT 10.010 -20.000 10.460 -19.920 ;
        RECT 8.160 -20.240 10.460 -20.000 ;
        RECT 8.160 -20.340 8.610 -20.240 ;
        RECT 10.010 -20.340 10.460 -20.240 ;
        RECT 11.410 -20.000 11.860 -19.890 ;
        RECT 13.260 -20.000 13.710 -19.890 ;
        RECT 11.410 -20.240 13.710 -20.000 ;
        RECT 11.410 -20.310 11.860 -20.240 ;
        RECT 5.420 -20.820 6.970 -20.600 ;
        RECT 5.420 -21.210 5.920 -20.820 ;
        RECT 6.520 -20.870 6.970 -20.820 ;
        RECT 7.350 -20.870 7.780 -20.810 ;
        RECT 8.160 -20.820 9.710 -20.600 ;
        RECT 12.460 -20.670 12.870 -20.240 ;
        RECT 13.260 -20.340 13.710 -20.240 ;
        RECT 14.920 -20.000 15.370 -19.890 ;
        RECT 16.770 -20.000 17.220 -19.890 ;
        RECT 14.920 -20.240 17.220 -20.000 ;
        RECT 14.920 -20.340 15.370 -20.240 ;
        RECT 15.760 -20.670 16.170 -20.240 ;
        RECT 16.770 -20.310 17.220 -20.240 ;
        RECT 18.170 -20.000 18.620 -19.920 ;
        RECT 19.220 -20.000 19.630 -19.560 ;
        RECT 20.020 -20.000 20.470 -19.890 ;
        RECT 18.170 -20.240 20.470 -20.000 ;
        RECT 18.170 -20.340 18.620 -20.240 ;
        RECT 20.020 -20.340 20.470 -20.240 ;
        RECT 21.660 -20.000 22.110 -19.890 ;
        RECT 22.500 -20.000 22.910 -19.560 ;
        RECT 25.680 -19.830 26.130 -19.550 ;
        RECT 29.500 -19.830 29.950 -19.550 ;
        RECT 39.180 -19.550 40.710 -19.340 ;
        RECT 41.090 -19.430 41.540 -19.340 ;
        RECT 41.920 -19.550 43.450 -19.340 ;
        RECT 23.510 -20.000 23.960 -19.920 ;
        RECT 21.660 -20.240 23.960 -20.000 ;
        RECT 21.660 -20.340 22.110 -20.240 ;
        RECT 23.510 -20.340 23.960 -20.240 ;
        RECT 24.910 -20.000 25.360 -19.890 ;
        RECT 26.760 -20.000 27.210 -19.890 ;
        RECT 24.910 -20.240 27.210 -20.000 ;
        RECT 24.910 -20.310 25.360 -20.240 ;
        RECT 8.160 -20.870 8.610 -20.820 ;
        RECT 6.520 -21.160 8.610 -20.870 ;
        RECT 6.520 -21.210 6.970 -21.160 ;
        RECT 1.420 -21.790 1.870 -21.690 ;
        RECT 2.260 -21.790 2.670 -21.360 ;
        RECT 5.420 -21.430 6.970 -21.210 ;
        RECT 7.350 -21.220 7.780 -21.160 ;
        RECT 8.160 -21.210 8.610 -21.160 ;
        RECT 9.210 -21.210 9.710 -20.820 ;
        RECT 8.160 -21.430 9.710 -21.210 ;
        RECT 18.920 -20.820 20.470 -20.600 ;
        RECT 18.920 -21.210 19.420 -20.820 ;
        RECT 20.020 -20.870 20.470 -20.820 ;
        RECT 20.850 -20.870 21.280 -20.810 ;
        RECT 21.660 -20.820 23.210 -20.600 ;
        RECT 25.960 -20.670 26.370 -20.240 ;
        RECT 26.760 -20.340 27.210 -20.240 ;
        RECT 28.420 -20.000 28.870 -19.890 ;
        RECT 30.270 -20.000 30.720 -19.890 ;
        RECT 28.420 -20.240 30.720 -20.000 ;
        RECT 28.420 -20.340 28.870 -20.240 ;
        RECT 29.260 -20.670 29.670 -20.240 ;
        RECT 30.270 -20.310 30.720 -20.240 ;
        RECT 31.670 -20.000 32.120 -19.920 ;
        RECT 32.720 -20.000 33.130 -19.560 ;
        RECT 33.520 -20.000 33.970 -19.890 ;
        RECT 31.670 -20.240 33.970 -20.000 ;
        RECT 31.670 -20.340 32.120 -20.240 ;
        RECT 33.520 -20.340 33.970 -20.240 ;
        RECT 35.160 -20.000 35.610 -19.890 ;
        RECT 36.000 -20.000 36.410 -19.560 ;
        RECT 39.180 -19.830 39.630 -19.550 ;
        RECT 43.000 -19.830 43.450 -19.550 ;
        RECT 52.680 -19.550 54.210 -19.340 ;
        RECT 54.590 -19.430 55.040 -19.340 ;
        RECT 55.420 -19.550 56.950 -19.340 ;
        RECT 37.010 -20.000 37.460 -19.920 ;
        RECT 35.160 -20.240 37.460 -20.000 ;
        RECT 35.160 -20.340 35.610 -20.240 ;
        RECT 37.010 -20.340 37.460 -20.240 ;
        RECT 38.410 -20.000 38.860 -19.890 ;
        RECT 40.260 -20.000 40.710 -19.890 ;
        RECT 38.410 -20.240 40.710 -20.000 ;
        RECT 38.410 -20.310 38.860 -20.240 ;
        RECT 21.660 -20.870 22.110 -20.820 ;
        RECT 20.020 -21.160 22.110 -20.870 ;
        RECT 20.020 -21.210 20.470 -21.160 ;
        RECT 3.270 -21.790 3.720 -21.720 ;
        RECT 1.420 -22.030 3.720 -21.790 ;
        RECT 1.420 -22.140 1.870 -22.030 ;
        RECT 3.270 -22.140 3.720 -22.030 ;
        RECT 4.670 -21.790 5.120 -21.690 ;
        RECT 6.520 -21.790 6.970 -21.690 ;
        RECT 4.670 -22.030 6.970 -21.790 ;
        RECT 4.670 -22.110 5.120 -22.030 ;
        RECT 5.720 -22.470 6.130 -22.030 ;
        RECT 6.520 -22.140 6.970 -22.030 ;
        RECT 8.160 -21.790 8.610 -21.690 ;
        RECT 10.010 -21.790 10.460 -21.690 ;
        RECT 8.160 -22.030 10.460 -21.790 ;
        RECT 8.160 -22.140 8.610 -22.030 ;
        RECT 9.000 -22.470 9.410 -22.030 ;
        RECT 10.010 -22.110 10.460 -22.030 ;
        RECT 11.410 -21.790 11.860 -21.720 ;
        RECT 12.460 -21.790 12.870 -21.360 ;
        RECT 13.260 -21.790 13.710 -21.690 ;
        RECT 11.410 -22.030 13.710 -21.790 ;
        RECT 11.410 -22.140 11.860 -22.030 ;
        RECT 13.260 -22.140 13.710 -22.030 ;
        RECT 14.920 -21.790 15.370 -21.690 ;
        RECT 15.760 -21.790 16.170 -21.360 ;
        RECT 18.920 -21.430 20.470 -21.210 ;
        RECT 20.850 -21.220 21.280 -21.160 ;
        RECT 21.660 -21.210 22.110 -21.160 ;
        RECT 22.710 -21.210 23.210 -20.820 ;
        RECT 21.660 -21.430 23.210 -21.210 ;
        RECT 32.420 -20.820 33.970 -20.600 ;
        RECT 32.420 -21.210 32.920 -20.820 ;
        RECT 33.520 -20.870 33.970 -20.820 ;
        RECT 34.350 -20.870 34.780 -20.810 ;
        RECT 35.160 -20.820 36.710 -20.600 ;
        RECT 39.460 -20.670 39.870 -20.240 ;
        RECT 40.260 -20.340 40.710 -20.240 ;
        RECT 41.920 -20.000 42.370 -19.890 ;
        RECT 43.770 -20.000 44.220 -19.890 ;
        RECT 41.920 -20.240 44.220 -20.000 ;
        RECT 41.920 -20.340 42.370 -20.240 ;
        RECT 42.760 -20.670 43.170 -20.240 ;
        RECT 43.770 -20.310 44.220 -20.240 ;
        RECT 45.170 -20.000 45.620 -19.920 ;
        RECT 46.220 -20.000 46.630 -19.560 ;
        RECT 47.020 -20.000 47.470 -19.890 ;
        RECT 45.170 -20.240 47.470 -20.000 ;
        RECT 45.170 -20.340 45.620 -20.240 ;
        RECT 47.020 -20.340 47.470 -20.240 ;
        RECT 48.660 -20.000 49.110 -19.890 ;
        RECT 49.500 -20.000 49.910 -19.560 ;
        RECT 52.680 -19.830 53.130 -19.550 ;
        RECT 56.500 -19.830 56.950 -19.550 ;
        RECT 66.180 -19.550 67.710 -19.340 ;
        RECT 68.090 -19.430 68.540 -19.340 ;
        RECT 68.920 -19.550 70.450 -19.340 ;
        RECT 50.510 -20.000 50.960 -19.920 ;
        RECT 48.660 -20.240 50.960 -20.000 ;
        RECT 48.660 -20.340 49.110 -20.240 ;
        RECT 50.510 -20.340 50.960 -20.240 ;
        RECT 51.910 -20.000 52.360 -19.890 ;
        RECT 53.760 -20.000 54.210 -19.890 ;
        RECT 51.910 -20.240 54.210 -20.000 ;
        RECT 51.910 -20.310 52.360 -20.240 ;
        RECT 35.160 -20.870 35.610 -20.820 ;
        RECT 33.520 -21.160 35.610 -20.870 ;
        RECT 33.520 -21.210 33.970 -21.160 ;
        RECT 16.770 -21.790 17.220 -21.720 ;
        RECT 14.920 -22.030 17.220 -21.790 ;
        RECT 14.920 -22.140 15.370 -22.030 ;
        RECT 16.770 -22.140 17.220 -22.030 ;
        RECT 18.170 -21.790 18.620 -21.690 ;
        RECT 20.020 -21.790 20.470 -21.690 ;
        RECT 18.170 -22.030 20.470 -21.790 ;
        RECT 18.170 -22.110 18.620 -22.030 ;
        RECT 12.180 -22.480 12.630 -22.200 ;
        RECT 16.000 -22.480 16.450 -22.200 ;
        RECT 19.220 -22.470 19.630 -22.030 ;
        RECT 20.020 -22.140 20.470 -22.030 ;
        RECT 21.660 -21.790 22.110 -21.690 ;
        RECT 23.510 -21.790 23.960 -21.690 ;
        RECT 21.660 -22.030 23.960 -21.790 ;
        RECT 21.660 -22.140 22.110 -22.030 ;
        RECT 22.500 -22.470 22.910 -22.030 ;
        RECT 23.510 -22.110 23.960 -22.030 ;
        RECT 24.910 -21.790 25.360 -21.720 ;
        RECT 25.960 -21.790 26.370 -21.360 ;
        RECT 26.760 -21.790 27.210 -21.690 ;
        RECT 24.910 -22.030 27.210 -21.790 ;
        RECT 24.910 -22.140 25.360 -22.030 ;
        RECT 26.760 -22.140 27.210 -22.030 ;
        RECT 28.420 -21.790 28.870 -21.690 ;
        RECT 29.260 -21.790 29.670 -21.360 ;
        RECT 32.420 -21.430 33.970 -21.210 ;
        RECT 34.350 -21.220 34.780 -21.160 ;
        RECT 35.160 -21.210 35.610 -21.160 ;
        RECT 36.210 -21.210 36.710 -20.820 ;
        RECT 35.160 -21.430 36.710 -21.210 ;
        RECT 45.920 -20.820 47.470 -20.600 ;
        RECT 45.920 -21.210 46.420 -20.820 ;
        RECT 47.020 -20.870 47.470 -20.820 ;
        RECT 47.850 -20.870 48.280 -20.810 ;
        RECT 48.660 -20.820 50.210 -20.600 ;
        RECT 52.960 -20.670 53.370 -20.240 ;
        RECT 53.760 -20.340 54.210 -20.240 ;
        RECT 55.420 -20.000 55.870 -19.890 ;
        RECT 57.270 -20.000 57.720 -19.890 ;
        RECT 55.420 -20.240 57.720 -20.000 ;
        RECT 55.420 -20.340 55.870 -20.240 ;
        RECT 56.260 -20.670 56.670 -20.240 ;
        RECT 57.270 -20.310 57.720 -20.240 ;
        RECT 58.670 -20.000 59.120 -19.920 ;
        RECT 59.720 -20.000 60.130 -19.560 ;
        RECT 60.520 -20.000 60.970 -19.890 ;
        RECT 58.670 -20.240 60.970 -20.000 ;
        RECT 58.670 -20.340 59.120 -20.240 ;
        RECT 60.520 -20.340 60.970 -20.240 ;
        RECT 62.160 -20.000 62.610 -19.890 ;
        RECT 63.000 -20.000 63.410 -19.560 ;
        RECT 66.180 -19.830 66.630 -19.550 ;
        RECT 70.000 -19.830 70.450 -19.550 ;
        RECT 79.680 -19.550 81.210 -19.340 ;
        RECT 81.590 -19.430 82.040 -19.340 ;
        RECT 82.420 -19.550 83.950 -19.340 ;
        RECT 64.010 -20.000 64.460 -19.920 ;
        RECT 62.160 -20.240 64.460 -20.000 ;
        RECT 62.160 -20.340 62.610 -20.240 ;
        RECT 64.010 -20.340 64.460 -20.240 ;
        RECT 65.410 -20.000 65.860 -19.890 ;
        RECT 67.260 -20.000 67.710 -19.890 ;
        RECT 65.410 -20.240 67.710 -20.000 ;
        RECT 65.410 -20.310 65.860 -20.240 ;
        RECT 48.660 -20.870 49.110 -20.820 ;
        RECT 47.020 -21.160 49.110 -20.870 ;
        RECT 47.020 -21.210 47.470 -21.160 ;
        RECT 30.270 -21.790 30.720 -21.720 ;
        RECT 28.420 -22.030 30.720 -21.790 ;
        RECT 28.420 -22.140 28.870 -22.030 ;
        RECT 30.270 -22.140 30.720 -22.030 ;
        RECT 31.670 -21.790 32.120 -21.690 ;
        RECT 33.520 -21.790 33.970 -21.690 ;
        RECT 31.670 -22.030 33.970 -21.790 ;
        RECT 31.670 -22.110 32.120 -22.030 ;
        RECT 12.180 -22.690 13.710 -22.480 ;
        RECT 14.090 -22.690 14.540 -22.600 ;
        RECT 14.920 -22.690 16.450 -22.480 ;
        RECT 25.680 -22.480 26.130 -22.200 ;
        RECT 29.500 -22.480 29.950 -22.200 ;
        RECT 32.720 -22.470 33.130 -22.030 ;
        RECT 33.520 -22.140 33.970 -22.030 ;
        RECT 35.160 -21.790 35.610 -21.690 ;
        RECT 37.010 -21.790 37.460 -21.690 ;
        RECT 35.160 -22.030 37.460 -21.790 ;
        RECT 35.160 -22.140 35.610 -22.030 ;
        RECT 36.000 -22.470 36.410 -22.030 ;
        RECT 37.010 -22.110 37.460 -22.030 ;
        RECT 38.410 -21.790 38.860 -21.720 ;
        RECT 39.460 -21.790 39.870 -21.360 ;
        RECT 40.260 -21.790 40.710 -21.690 ;
        RECT 38.410 -22.030 40.710 -21.790 ;
        RECT 38.410 -22.140 38.860 -22.030 ;
        RECT 40.260 -22.140 40.710 -22.030 ;
        RECT 41.920 -21.790 42.370 -21.690 ;
        RECT 42.760 -21.790 43.170 -21.360 ;
        RECT 45.920 -21.430 47.470 -21.210 ;
        RECT 47.850 -21.220 48.280 -21.160 ;
        RECT 48.660 -21.210 49.110 -21.160 ;
        RECT 49.710 -21.210 50.210 -20.820 ;
        RECT 48.660 -21.430 50.210 -21.210 ;
        RECT 59.420 -20.820 60.970 -20.600 ;
        RECT 59.420 -21.210 59.920 -20.820 ;
        RECT 60.520 -20.870 60.970 -20.820 ;
        RECT 61.350 -20.870 61.780 -20.810 ;
        RECT 62.160 -20.820 63.710 -20.600 ;
        RECT 66.460 -20.670 66.870 -20.240 ;
        RECT 67.260 -20.340 67.710 -20.240 ;
        RECT 68.920 -20.000 69.370 -19.890 ;
        RECT 70.770 -20.000 71.220 -19.890 ;
        RECT 68.920 -20.240 71.220 -20.000 ;
        RECT 68.920 -20.340 69.370 -20.240 ;
        RECT 69.760 -20.670 70.170 -20.240 ;
        RECT 70.770 -20.310 71.220 -20.240 ;
        RECT 72.170 -20.000 72.620 -19.920 ;
        RECT 73.220 -20.000 73.630 -19.560 ;
        RECT 74.020 -20.000 74.470 -19.890 ;
        RECT 72.170 -20.240 74.470 -20.000 ;
        RECT 72.170 -20.340 72.620 -20.240 ;
        RECT 74.020 -20.340 74.470 -20.240 ;
        RECT 75.660 -20.000 76.110 -19.890 ;
        RECT 76.500 -20.000 76.910 -19.560 ;
        RECT 79.680 -19.830 80.130 -19.550 ;
        RECT 83.500 -19.830 83.950 -19.550 ;
        RECT 93.180 -19.550 94.710 -19.340 ;
        RECT 95.090 -19.430 95.540 -19.340 ;
        RECT 95.920 -19.550 97.450 -19.340 ;
        RECT 77.510 -20.000 77.960 -19.920 ;
        RECT 75.660 -20.240 77.960 -20.000 ;
        RECT 75.660 -20.340 76.110 -20.240 ;
        RECT 77.510 -20.340 77.960 -20.240 ;
        RECT 78.910 -20.000 79.360 -19.890 ;
        RECT 80.760 -20.000 81.210 -19.890 ;
        RECT 78.910 -20.240 81.210 -20.000 ;
        RECT 78.910 -20.310 79.360 -20.240 ;
        RECT 62.160 -20.870 62.610 -20.820 ;
        RECT 60.520 -21.160 62.610 -20.870 ;
        RECT 60.520 -21.210 60.970 -21.160 ;
        RECT 43.770 -21.790 44.220 -21.720 ;
        RECT 41.920 -22.030 44.220 -21.790 ;
        RECT 41.920 -22.140 42.370 -22.030 ;
        RECT 43.770 -22.140 44.220 -22.030 ;
        RECT 45.170 -21.790 45.620 -21.690 ;
        RECT 47.020 -21.790 47.470 -21.690 ;
        RECT 45.170 -22.030 47.470 -21.790 ;
        RECT 45.170 -22.110 45.620 -22.030 ;
        RECT 25.680 -22.690 27.210 -22.480 ;
        RECT 27.590 -22.690 28.040 -22.600 ;
        RECT 28.420 -22.690 29.950 -22.480 ;
        RECT 39.180 -22.480 39.630 -22.200 ;
        RECT 43.000 -22.480 43.450 -22.200 ;
        RECT 46.220 -22.470 46.630 -22.030 ;
        RECT 47.020 -22.140 47.470 -22.030 ;
        RECT 48.660 -21.790 49.110 -21.690 ;
        RECT 50.510 -21.790 50.960 -21.690 ;
        RECT 48.660 -22.030 50.960 -21.790 ;
        RECT 48.660 -22.140 49.110 -22.030 ;
        RECT 49.500 -22.470 49.910 -22.030 ;
        RECT 50.510 -22.110 50.960 -22.030 ;
        RECT 51.910 -21.790 52.360 -21.720 ;
        RECT 52.960 -21.790 53.370 -21.360 ;
        RECT 53.760 -21.790 54.210 -21.690 ;
        RECT 51.910 -22.030 54.210 -21.790 ;
        RECT 51.910 -22.140 52.360 -22.030 ;
        RECT 53.760 -22.140 54.210 -22.030 ;
        RECT 55.420 -21.790 55.870 -21.690 ;
        RECT 56.260 -21.790 56.670 -21.360 ;
        RECT 59.420 -21.430 60.970 -21.210 ;
        RECT 61.350 -21.220 61.780 -21.160 ;
        RECT 62.160 -21.210 62.610 -21.160 ;
        RECT 63.210 -21.210 63.710 -20.820 ;
        RECT 62.160 -21.430 63.710 -21.210 ;
        RECT 72.920 -20.820 74.470 -20.600 ;
        RECT 72.920 -21.210 73.420 -20.820 ;
        RECT 74.020 -20.870 74.470 -20.820 ;
        RECT 74.850 -20.870 75.280 -20.810 ;
        RECT 75.660 -20.820 77.210 -20.600 ;
        RECT 79.960 -20.670 80.370 -20.240 ;
        RECT 80.760 -20.340 81.210 -20.240 ;
        RECT 82.420 -20.000 82.870 -19.890 ;
        RECT 84.270 -20.000 84.720 -19.890 ;
        RECT 82.420 -20.240 84.720 -20.000 ;
        RECT 82.420 -20.340 82.870 -20.240 ;
        RECT 83.260 -20.670 83.670 -20.240 ;
        RECT 84.270 -20.310 84.720 -20.240 ;
        RECT 85.670 -20.000 86.120 -19.920 ;
        RECT 86.720 -20.000 87.130 -19.560 ;
        RECT 87.520 -20.000 87.970 -19.890 ;
        RECT 85.670 -20.240 87.970 -20.000 ;
        RECT 85.670 -20.340 86.120 -20.240 ;
        RECT 87.520 -20.340 87.970 -20.240 ;
        RECT 89.160 -20.000 89.610 -19.890 ;
        RECT 90.000 -20.000 90.410 -19.560 ;
        RECT 93.180 -19.830 93.630 -19.550 ;
        RECT 97.000 -19.830 97.450 -19.550 ;
        RECT 106.680 -19.550 108.210 -19.340 ;
        RECT 108.590 -19.430 109.040 -19.340 ;
        RECT 109.420 -19.550 110.950 -19.340 ;
        RECT 91.010 -20.000 91.460 -19.920 ;
        RECT 89.160 -20.240 91.460 -20.000 ;
        RECT 89.160 -20.340 89.610 -20.240 ;
        RECT 91.010 -20.340 91.460 -20.240 ;
        RECT 92.410 -20.000 92.860 -19.890 ;
        RECT 94.260 -20.000 94.710 -19.890 ;
        RECT 92.410 -20.240 94.710 -20.000 ;
        RECT 92.410 -20.310 92.860 -20.240 ;
        RECT 75.660 -20.870 76.110 -20.820 ;
        RECT 74.020 -21.160 76.110 -20.870 ;
        RECT 74.020 -21.210 74.470 -21.160 ;
        RECT 57.270 -21.790 57.720 -21.720 ;
        RECT 55.420 -22.030 57.720 -21.790 ;
        RECT 55.420 -22.140 55.870 -22.030 ;
        RECT 57.270 -22.140 57.720 -22.030 ;
        RECT 58.670 -21.790 59.120 -21.690 ;
        RECT 60.520 -21.790 60.970 -21.690 ;
        RECT 58.670 -22.030 60.970 -21.790 ;
        RECT 58.670 -22.110 59.120 -22.030 ;
        RECT 39.180 -22.690 40.710 -22.480 ;
        RECT 41.090 -22.690 41.540 -22.600 ;
        RECT 41.920 -22.690 43.450 -22.480 ;
        RECT 52.680 -22.480 53.130 -22.200 ;
        RECT 56.500 -22.480 56.950 -22.200 ;
        RECT 59.720 -22.470 60.130 -22.030 ;
        RECT 60.520 -22.140 60.970 -22.030 ;
        RECT 62.160 -21.790 62.610 -21.690 ;
        RECT 64.010 -21.790 64.460 -21.690 ;
        RECT 62.160 -22.030 64.460 -21.790 ;
        RECT 62.160 -22.140 62.610 -22.030 ;
        RECT 63.000 -22.470 63.410 -22.030 ;
        RECT 64.010 -22.110 64.460 -22.030 ;
        RECT 65.410 -21.790 65.860 -21.720 ;
        RECT 66.460 -21.790 66.870 -21.360 ;
        RECT 67.260 -21.790 67.710 -21.690 ;
        RECT 65.410 -22.030 67.710 -21.790 ;
        RECT 65.410 -22.140 65.860 -22.030 ;
        RECT 67.260 -22.140 67.710 -22.030 ;
        RECT 68.920 -21.790 69.370 -21.690 ;
        RECT 69.760 -21.790 70.170 -21.360 ;
        RECT 72.920 -21.430 74.470 -21.210 ;
        RECT 74.850 -21.220 75.280 -21.160 ;
        RECT 75.660 -21.210 76.110 -21.160 ;
        RECT 76.710 -21.210 77.210 -20.820 ;
        RECT 75.660 -21.430 77.210 -21.210 ;
        RECT 86.420 -20.820 87.970 -20.600 ;
        RECT 86.420 -21.210 86.920 -20.820 ;
        RECT 87.520 -20.870 87.970 -20.820 ;
        RECT 88.350 -20.870 88.780 -20.810 ;
        RECT 89.160 -20.820 90.710 -20.600 ;
        RECT 93.460 -20.670 93.870 -20.240 ;
        RECT 94.260 -20.340 94.710 -20.240 ;
        RECT 95.920 -20.000 96.370 -19.890 ;
        RECT 97.770 -20.000 98.220 -19.890 ;
        RECT 95.920 -20.240 98.220 -20.000 ;
        RECT 95.920 -20.340 96.370 -20.240 ;
        RECT 96.760 -20.670 97.170 -20.240 ;
        RECT 97.770 -20.310 98.220 -20.240 ;
        RECT 99.170 -20.000 99.620 -19.920 ;
        RECT 100.220 -20.000 100.630 -19.560 ;
        RECT 101.020 -20.000 101.470 -19.890 ;
        RECT 99.170 -20.240 101.470 -20.000 ;
        RECT 99.170 -20.340 99.620 -20.240 ;
        RECT 101.020 -20.340 101.470 -20.240 ;
        RECT 102.660 -20.000 103.110 -19.890 ;
        RECT 103.500 -20.000 103.910 -19.560 ;
        RECT 106.680 -19.830 107.130 -19.550 ;
        RECT 110.500 -19.830 110.950 -19.550 ;
        RECT 120.180 -19.550 121.710 -19.340 ;
        RECT 122.090 -19.430 122.540 -19.340 ;
        RECT 122.920 -19.550 124.450 -19.340 ;
        RECT 104.510 -20.000 104.960 -19.920 ;
        RECT 102.660 -20.240 104.960 -20.000 ;
        RECT 102.660 -20.340 103.110 -20.240 ;
        RECT 104.510 -20.340 104.960 -20.240 ;
        RECT 105.910 -20.000 106.360 -19.890 ;
        RECT 107.760 -20.000 108.210 -19.890 ;
        RECT 105.910 -20.240 108.210 -20.000 ;
        RECT 105.910 -20.310 106.360 -20.240 ;
        RECT 89.160 -20.870 89.610 -20.820 ;
        RECT 87.520 -21.160 89.610 -20.870 ;
        RECT 87.520 -21.210 87.970 -21.160 ;
        RECT 70.770 -21.790 71.220 -21.720 ;
        RECT 68.920 -22.030 71.220 -21.790 ;
        RECT 68.920 -22.140 69.370 -22.030 ;
        RECT 70.770 -22.140 71.220 -22.030 ;
        RECT 72.170 -21.790 72.620 -21.690 ;
        RECT 74.020 -21.790 74.470 -21.690 ;
        RECT 72.170 -22.030 74.470 -21.790 ;
        RECT 72.170 -22.110 72.620 -22.030 ;
        RECT 52.680 -22.690 54.210 -22.480 ;
        RECT 54.590 -22.690 55.040 -22.600 ;
        RECT 55.420 -22.690 56.950 -22.480 ;
        RECT 66.180 -22.480 66.630 -22.200 ;
        RECT 70.000 -22.480 70.450 -22.200 ;
        RECT 73.220 -22.470 73.630 -22.030 ;
        RECT 74.020 -22.140 74.470 -22.030 ;
        RECT 75.660 -21.790 76.110 -21.690 ;
        RECT 77.510 -21.790 77.960 -21.690 ;
        RECT 75.660 -22.030 77.960 -21.790 ;
        RECT 75.660 -22.140 76.110 -22.030 ;
        RECT 76.500 -22.470 76.910 -22.030 ;
        RECT 77.510 -22.110 77.960 -22.030 ;
        RECT 78.910 -21.790 79.360 -21.720 ;
        RECT 79.960 -21.790 80.370 -21.360 ;
        RECT 80.760 -21.790 81.210 -21.690 ;
        RECT 78.910 -22.030 81.210 -21.790 ;
        RECT 78.910 -22.140 79.360 -22.030 ;
        RECT 80.760 -22.140 81.210 -22.030 ;
        RECT 82.420 -21.790 82.870 -21.690 ;
        RECT 83.260 -21.790 83.670 -21.360 ;
        RECT 86.420 -21.430 87.970 -21.210 ;
        RECT 88.350 -21.220 88.780 -21.160 ;
        RECT 89.160 -21.210 89.610 -21.160 ;
        RECT 90.210 -21.210 90.710 -20.820 ;
        RECT 89.160 -21.430 90.710 -21.210 ;
        RECT 99.920 -20.820 101.470 -20.600 ;
        RECT 99.920 -21.210 100.420 -20.820 ;
        RECT 101.020 -20.870 101.470 -20.820 ;
        RECT 101.850 -20.870 102.280 -20.810 ;
        RECT 102.660 -20.820 104.210 -20.600 ;
        RECT 106.960 -20.670 107.370 -20.240 ;
        RECT 107.760 -20.340 108.210 -20.240 ;
        RECT 109.420 -20.000 109.870 -19.890 ;
        RECT 111.270 -20.000 111.720 -19.890 ;
        RECT 109.420 -20.240 111.720 -20.000 ;
        RECT 109.420 -20.340 109.870 -20.240 ;
        RECT 110.260 -20.670 110.670 -20.240 ;
        RECT 111.270 -20.310 111.720 -20.240 ;
        RECT 112.670 -20.000 113.120 -19.920 ;
        RECT 113.720 -20.000 114.130 -19.560 ;
        RECT 114.520 -20.000 114.970 -19.890 ;
        RECT 112.670 -20.240 114.970 -20.000 ;
        RECT 112.670 -20.340 113.120 -20.240 ;
        RECT 114.520 -20.340 114.970 -20.240 ;
        RECT 116.160 -20.000 116.610 -19.890 ;
        RECT 117.000 -20.000 117.410 -19.560 ;
        RECT 120.180 -19.830 120.630 -19.550 ;
        RECT 124.000 -19.830 124.450 -19.550 ;
        RECT 133.680 -19.550 135.210 -19.340 ;
        RECT 135.590 -19.430 136.040 -19.340 ;
        RECT 136.420 -19.550 137.950 -19.340 ;
        RECT 118.010 -20.000 118.460 -19.920 ;
        RECT 116.160 -20.240 118.460 -20.000 ;
        RECT 116.160 -20.340 116.610 -20.240 ;
        RECT 118.010 -20.340 118.460 -20.240 ;
        RECT 119.410 -20.000 119.860 -19.890 ;
        RECT 121.260 -20.000 121.710 -19.890 ;
        RECT 119.410 -20.240 121.710 -20.000 ;
        RECT 119.410 -20.310 119.860 -20.240 ;
        RECT 102.660 -20.870 103.110 -20.820 ;
        RECT 101.020 -21.160 103.110 -20.870 ;
        RECT 101.020 -21.210 101.470 -21.160 ;
        RECT 84.270 -21.790 84.720 -21.720 ;
        RECT 82.420 -22.030 84.720 -21.790 ;
        RECT 82.420 -22.140 82.870 -22.030 ;
        RECT 84.270 -22.140 84.720 -22.030 ;
        RECT 85.670 -21.790 86.120 -21.690 ;
        RECT 87.520 -21.790 87.970 -21.690 ;
        RECT 85.670 -22.030 87.970 -21.790 ;
        RECT 85.670 -22.110 86.120 -22.030 ;
        RECT 66.180 -22.690 67.710 -22.480 ;
        RECT 68.090 -22.690 68.540 -22.600 ;
        RECT 68.920 -22.690 70.450 -22.480 ;
        RECT 79.680 -22.480 80.130 -22.200 ;
        RECT 83.500 -22.480 83.950 -22.200 ;
        RECT 86.720 -22.470 87.130 -22.030 ;
        RECT 87.520 -22.140 87.970 -22.030 ;
        RECT 89.160 -21.790 89.610 -21.690 ;
        RECT 91.010 -21.790 91.460 -21.690 ;
        RECT 89.160 -22.030 91.460 -21.790 ;
        RECT 89.160 -22.140 89.610 -22.030 ;
        RECT 90.000 -22.470 90.410 -22.030 ;
        RECT 91.010 -22.110 91.460 -22.030 ;
        RECT 92.410 -21.790 92.860 -21.720 ;
        RECT 93.460 -21.790 93.870 -21.360 ;
        RECT 94.260 -21.790 94.710 -21.690 ;
        RECT 92.410 -22.030 94.710 -21.790 ;
        RECT 92.410 -22.140 92.860 -22.030 ;
        RECT 94.260 -22.140 94.710 -22.030 ;
        RECT 95.920 -21.790 96.370 -21.690 ;
        RECT 96.760 -21.790 97.170 -21.360 ;
        RECT 99.920 -21.430 101.470 -21.210 ;
        RECT 101.850 -21.220 102.280 -21.160 ;
        RECT 102.660 -21.210 103.110 -21.160 ;
        RECT 103.710 -21.210 104.210 -20.820 ;
        RECT 102.660 -21.430 104.210 -21.210 ;
        RECT 113.420 -20.820 114.970 -20.600 ;
        RECT 113.420 -21.210 113.920 -20.820 ;
        RECT 114.520 -20.870 114.970 -20.820 ;
        RECT 115.350 -20.870 115.780 -20.810 ;
        RECT 116.160 -20.820 117.710 -20.600 ;
        RECT 120.460 -20.670 120.870 -20.240 ;
        RECT 121.260 -20.340 121.710 -20.240 ;
        RECT 122.920 -20.000 123.370 -19.890 ;
        RECT 124.770 -20.000 125.220 -19.890 ;
        RECT 122.920 -20.240 125.220 -20.000 ;
        RECT 122.920 -20.340 123.370 -20.240 ;
        RECT 123.760 -20.670 124.170 -20.240 ;
        RECT 124.770 -20.310 125.220 -20.240 ;
        RECT 126.170 -20.000 126.620 -19.920 ;
        RECT 127.220 -20.000 127.630 -19.560 ;
        RECT 128.020 -20.000 128.470 -19.890 ;
        RECT 126.170 -20.240 128.470 -20.000 ;
        RECT 126.170 -20.340 126.620 -20.240 ;
        RECT 128.020 -20.340 128.470 -20.240 ;
        RECT 129.660 -20.000 130.110 -19.890 ;
        RECT 130.500 -20.000 130.910 -19.560 ;
        RECT 133.680 -19.830 134.130 -19.550 ;
        RECT 137.500 -19.830 137.950 -19.550 ;
        RECT 147.180 -19.550 148.710 -19.340 ;
        RECT 149.090 -19.430 149.540 -19.340 ;
        RECT 149.920 -19.550 151.450 -19.340 ;
        RECT 131.510 -20.000 131.960 -19.920 ;
        RECT 129.660 -20.240 131.960 -20.000 ;
        RECT 129.660 -20.340 130.110 -20.240 ;
        RECT 131.510 -20.340 131.960 -20.240 ;
        RECT 132.910 -20.000 133.360 -19.890 ;
        RECT 134.760 -20.000 135.210 -19.890 ;
        RECT 132.910 -20.240 135.210 -20.000 ;
        RECT 132.910 -20.310 133.360 -20.240 ;
        RECT 116.160 -20.870 116.610 -20.820 ;
        RECT 114.520 -21.160 116.610 -20.870 ;
        RECT 114.520 -21.210 114.970 -21.160 ;
        RECT 97.770 -21.790 98.220 -21.720 ;
        RECT 95.920 -22.030 98.220 -21.790 ;
        RECT 95.920 -22.140 96.370 -22.030 ;
        RECT 97.770 -22.140 98.220 -22.030 ;
        RECT 99.170 -21.790 99.620 -21.690 ;
        RECT 101.020 -21.790 101.470 -21.690 ;
        RECT 99.170 -22.030 101.470 -21.790 ;
        RECT 99.170 -22.110 99.620 -22.030 ;
        RECT 79.680 -22.690 81.210 -22.480 ;
        RECT 81.590 -22.690 82.040 -22.600 ;
        RECT 82.420 -22.690 83.950 -22.480 ;
        RECT 93.180 -22.480 93.630 -22.200 ;
        RECT 97.000 -22.480 97.450 -22.200 ;
        RECT 100.220 -22.470 100.630 -22.030 ;
        RECT 101.020 -22.140 101.470 -22.030 ;
        RECT 102.660 -21.790 103.110 -21.690 ;
        RECT 104.510 -21.790 104.960 -21.690 ;
        RECT 102.660 -22.030 104.960 -21.790 ;
        RECT 102.660 -22.140 103.110 -22.030 ;
        RECT 103.500 -22.470 103.910 -22.030 ;
        RECT 104.510 -22.110 104.960 -22.030 ;
        RECT 105.910 -21.790 106.360 -21.720 ;
        RECT 106.960 -21.790 107.370 -21.360 ;
        RECT 107.760 -21.790 108.210 -21.690 ;
        RECT 105.910 -22.030 108.210 -21.790 ;
        RECT 105.910 -22.140 106.360 -22.030 ;
        RECT 107.760 -22.140 108.210 -22.030 ;
        RECT 109.420 -21.790 109.870 -21.690 ;
        RECT 110.260 -21.790 110.670 -21.360 ;
        RECT 113.420 -21.430 114.970 -21.210 ;
        RECT 115.350 -21.220 115.780 -21.160 ;
        RECT 116.160 -21.210 116.610 -21.160 ;
        RECT 117.210 -21.210 117.710 -20.820 ;
        RECT 116.160 -21.430 117.710 -21.210 ;
        RECT 126.920 -20.820 128.470 -20.600 ;
        RECT 126.920 -21.210 127.420 -20.820 ;
        RECT 128.020 -20.870 128.470 -20.820 ;
        RECT 128.850 -20.870 129.280 -20.810 ;
        RECT 129.660 -20.820 131.210 -20.600 ;
        RECT 133.960 -20.670 134.370 -20.240 ;
        RECT 134.760 -20.340 135.210 -20.240 ;
        RECT 136.420 -20.000 136.870 -19.890 ;
        RECT 138.270 -20.000 138.720 -19.890 ;
        RECT 136.420 -20.240 138.720 -20.000 ;
        RECT 136.420 -20.340 136.870 -20.240 ;
        RECT 137.260 -20.670 137.670 -20.240 ;
        RECT 138.270 -20.310 138.720 -20.240 ;
        RECT 139.670 -20.000 140.120 -19.920 ;
        RECT 140.720 -20.000 141.130 -19.560 ;
        RECT 141.520 -20.000 141.970 -19.890 ;
        RECT 139.670 -20.240 141.970 -20.000 ;
        RECT 139.670 -20.340 140.120 -20.240 ;
        RECT 141.520 -20.340 141.970 -20.240 ;
        RECT 143.160 -20.000 143.610 -19.890 ;
        RECT 144.000 -20.000 144.410 -19.560 ;
        RECT 147.180 -19.830 147.630 -19.550 ;
        RECT 151.000 -19.830 151.450 -19.550 ;
        RECT 160.680 -19.550 162.210 -19.340 ;
        RECT 162.590 -19.430 163.040 -19.340 ;
        RECT 163.420 -19.550 164.950 -19.340 ;
        RECT 145.010 -20.000 145.460 -19.920 ;
        RECT 143.160 -20.240 145.460 -20.000 ;
        RECT 143.160 -20.340 143.610 -20.240 ;
        RECT 145.010 -20.340 145.460 -20.240 ;
        RECT 146.410 -20.000 146.860 -19.890 ;
        RECT 148.260 -20.000 148.710 -19.890 ;
        RECT 146.410 -20.240 148.710 -20.000 ;
        RECT 146.410 -20.310 146.860 -20.240 ;
        RECT 129.660 -20.870 130.110 -20.820 ;
        RECT 128.020 -21.160 130.110 -20.870 ;
        RECT 128.020 -21.210 128.470 -21.160 ;
        RECT 111.270 -21.790 111.720 -21.720 ;
        RECT 109.420 -22.030 111.720 -21.790 ;
        RECT 109.420 -22.140 109.870 -22.030 ;
        RECT 111.270 -22.140 111.720 -22.030 ;
        RECT 112.670 -21.790 113.120 -21.690 ;
        RECT 114.520 -21.790 114.970 -21.690 ;
        RECT 112.670 -22.030 114.970 -21.790 ;
        RECT 112.670 -22.110 113.120 -22.030 ;
        RECT 93.180 -22.690 94.710 -22.480 ;
        RECT 95.090 -22.690 95.540 -22.600 ;
        RECT 95.920 -22.690 97.450 -22.480 ;
        RECT 106.680 -22.480 107.130 -22.200 ;
        RECT 110.500 -22.480 110.950 -22.200 ;
        RECT 113.720 -22.470 114.130 -22.030 ;
        RECT 114.520 -22.140 114.970 -22.030 ;
        RECT 116.160 -21.790 116.610 -21.690 ;
        RECT 118.010 -21.790 118.460 -21.690 ;
        RECT 116.160 -22.030 118.460 -21.790 ;
        RECT 116.160 -22.140 116.610 -22.030 ;
        RECT 117.000 -22.470 117.410 -22.030 ;
        RECT 118.010 -22.110 118.460 -22.030 ;
        RECT 119.410 -21.790 119.860 -21.720 ;
        RECT 120.460 -21.790 120.870 -21.360 ;
        RECT 121.260 -21.790 121.710 -21.690 ;
        RECT 119.410 -22.030 121.710 -21.790 ;
        RECT 119.410 -22.140 119.860 -22.030 ;
        RECT 121.260 -22.140 121.710 -22.030 ;
        RECT 122.920 -21.790 123.370 -21.690 ;
        RECT 123.760 -21.790 124.170 -21.360 ;
        RECT 126.920 -21.430 128.470 -21.210 ;
        RECT 128.850 -21.220 129.280 -21.160 ;
        RECT 129.660 -21.210 130.110 -21.160 ;
        RECT 130.710 -21.210 131.210 -20.820 ;
        RECT 129.660 -21.430 131.210 -21.210 ;
        RECT 140.420 -20.820 141.970 -20.600 ;
        RECT 140.420 -21.210 140.920 -20.820 ;
        RECT 141.520 -20.870 141.970 -20.820 ;
        RECT 142.350 -20.870 142.780 -20.810 ;
        RECT 143.160 -20.820 144.710 -20.600 ;
        RECT 147.460 -20.670 147.870 -20.240 ;
        RECT 148.260 -20.340 148.710 -20.240 ;
        RECT 149.920 -20.000 150.370 -19.890 ;
        RECT 151.770 -20.000 152.220 -19.890 ;
        RECT 149.920 -20.240 152.220 -20.000 ;
        RECT 149.920 -20.340 150.370 -20.240 ;
        RECT 150.760 -20.670 151.170 -20.240 ;
        RECT 151.770 -20.310 152.220 -20.240 ;
        RECT 153.170 -20.000 153.620 -19.920 ;
        RECT 154.220 -20.000 154.630 -19.560 ;
        RECT 155.020 -20.000 155.470 -19.890 ;
        RECT 153.170 -20.240 155.470 -20.000 ;
        RECT 153.170 -20.340 153.620 -20.240 ;
        RECT 155.020 -20.340 155.470 -20.240 ;
        RECT 156.660 -20.000 157.110 -19.890 ;
        RECT 157.500 -20.000 157.910 -19.560 ;
        RECT 160.680 -19.830 161.130 -19.550 ;
        RECT 164.500 -19.830 164.950 -19.550 ;
        RECT 174.180 -19.550 175.710 -19.340 ;
        RECT 176.090 -19.430 176.540 -19.340 ;
        RECT 176.920 -19.550 178.450 -19.340 ;
        RECT 158.510 -20.000 158.960 -19.920 ;
        RECT 156.660 -20.240 158.960 -20.000 ;
        RECT 156.660 -20.340 157.110 -20.240 ;
        RECT 158.510 -20.340 158.960 -20.240 ;
        RECT 159.910 -20.000 160.360 -19.890 ;
        RECT 161.760 -20.000 162.210 -19.890 ;
        RECT 159.910 -20.240 162.210 -20.000 ;
        RECT 159.910 -20.310 160.360 -20.240 ;
        RECT 143.160 -20.870 143.610 -20.820 ;
        RECT 141.520 -21.160 143.610 -20.870 ;
        RECT 141.520 -21.210 141.970 -21.160 ;
        RECT 124.770 -21.790 125.220 -21.720 ;
        RECT 122.920 -22.030 125.220 -21.790 ;
        RECT 122.920 -22.140 123.370 -22.030 ;
        RECT 124.770 -22.140 125.220 -22.030 ;
        RECT 126.170 -21.790 126.620 -21.690 ;
        RECT 128.020 -21.790 128.470 -21.690 ;
        RECT 126.170 -22.030 128.470 -21.790 ;
        RECT 126.170 -22.110 126.620 -22.030 ;
        RECT 106.680 -22.690 108.210 -22.480 ;
        RECT 108.590 -22.690 109.040 -22.600 ;
        RECT 109.420 -22.690 110.950 -22.480 ;
        RECT 120.180 -22.480 120.630 -22.200 ;
        RECT 124.000 -22.480 124.450 -22.200 ;
        RECT 127.220 -22.470 127.630 -22.030 ;
        RECT 128.020 -22.140 128.470 -22.030 ;
        RECT 129.660 -21.790 130.110 -21.690 ;
        RECT 131.510 -21.790 131.960 -21.690 ;
        RECT 129.660 -22.030 131.960 -21.790 ;
        RECT 129.660 -22.140 130.110 -22.030 ;
        RECT 130.500 -22.470 130.910 -22.030 ;
        RECT 131.510 -22.110 131.960 -22.030 ;
        RECT 132.910 -21.790 133.360 -21.720 ;
        RECT 133.960 -21.790 134.370 -21.360 ;
        RECT 134.760 -21.790 135.210 -21.690 ;
        RECT 132.910 -22.030 135.210 -21.790 ;
        RECT 132.910 -22.140 133.360 -22.030 ;
        RECT 134.760 -22.140 135.210 -22.030 ;
        RECT 136.420 -21.790 136.870 -21.690 ;
        RECT 137.260 -21.790 137.670 -21.360 ;
        RECT 140.420 -21.430 141.970 -21.210 ;
        RECT 142.350 -21.220 142.780 -21.160 ;
        RECT 143.160 -21.210 143.610 -21.160 ;
        RECT 144.210 -21.210 144.710 -20.820 ;
        RECT 143.160 -21.430 144.710 -21.210 ;
        RECT 153.920 -20.820 155.470 -20.600 ;
        RECT 153.920 -21.210 154.420 -20.820 ;
        RECT 155.020 -20.870 155.470 -20.820 ;
        RECT 155.850 -20.870 156.280 -20.810 ;
        RECT 156.660 -20.820 158.210 -20.600 ;
        RECT 160.960 -20.670 161.370 -20.240 ;
        RECT 161.760 -20.340 162.210 -20.240 ;
        RECT 163.420 -20.000 163.870 -19.890 ;
        RECT 165.270 -20.000 165.720 -19.890 ;
        RECT 163.420 -20.240 165.720 -20.000 ;
        RECT 163.420 -20.340 163.870 -20.240 ;
        RECT 164.260 -20.670 164.670 -20.240 ;
        RECT 165.270 -20.310 165.720 -20.240 ;
        RECT 166.670 -20.000 167.120 -19.920 ;
        RECT 167.720 -20.000 168.130 -19.560 ;
        RECT 168.520 -20.000 168.970 -19.890 ;
        RECT 166.670 -20.240 168.970 -20.000 ;
        RECT 166.670 -20.340 167.120 -20.240 ;
        RECT 168.520 -20.340 168.970 -20.240 ;
        RECT 170.160 -20.000 170.610 -19.890 ;
        RECT 171.000 -20.000 171.410 -19.560 ;
        RECT 174.180 -19.830 174.630 -19.550 ;
        RECT 178.000 -19.830 178.450 -19.550 ;
        RECT 187.680 -19.550 189.210 -19.340 ;
        RECT 189.590 -19.430 190.040 -19.340 ;
        RECT 190.420 -19.550 191.950 -19.340 ;
        RECT 172.010 -20.000 172.460 -19.920 ;
        RECT 170.160 -20.240 172.460 -20.000 ;
        RECT 170.160 -20.340 170.610 -20.240 ;
        RECT 172.010 -20.340 172.460 -20.240 ;
        RECT 173.410 -20.000 173.860 -19.890 ;
        RECT 175.260 -20.000 175.710 -19.890 ;
        RECT 173.410 -20.240 175.710 -20.000 ;
        RECT 173.410 -20.310 173.860 -20.240 ;
        RECT 156.660 -20.870 157.110 -20.820 ;
        RECT 155.020 -21.160 157.110 -20.870 ;
        RECT 155.020 -21.210 155.470 -21.160 ;
        RECT 138.270 -21.790 138.720 -21.720 ;
        RECT 136.420 -22.030 138.720 -21.790 ;
        RECT 136.420 -22.140 136.870 -22.030 ;
        RECT 138.270 -22.140 138.720 -22.030 ;
        RECT 139.670 -21.790 140.120 -21.690 ;
        RECT 141.520 -21.790 141.970 -21.690 ;
        RECT 139.670 -22.030 141.970 -21.790 ;
        RECT 139.670 -22.110 140.120 -22.030 ;
        RECT 120.180 -22.690 121.710 -22.480 ;
        RECT 122.090 -22.690 122.540 -22.600 ;
        RECT 122.920 -22.690 124.450 -22.480 ;
        RECT 133.680 -22.480 134.130 -22.200 ;
        RECT 137.500 -22.480 137.950 -22.200 ;
        RECT 140.720 -22.470 141.130 -22.030 ;
        RECT 141.520 -22.140 141.970 -22.030 ;
        RECT 143.160 -21.790 143.610 -21.690 ;
        RECT 145.010 -21.790 145.460 -21.690 ;
        RECT 143.160 -22.030 145.460 -21.790 ;
        RECT 143.160 -22.140 143.610 -22.030 ;
        RECT 144.000 -22.470 144.410 -22.030 ;
        RECT 145.010 -22.110 145.460 -22.030 ;
        RECT 146.410 -21.790 146.860 -21.720 ;
        RECT 147.460 -21.790 147.870 -21.360 ;
        RECT 148.260 -21.790 148.710 -21.690 ;
        RECT 146.410 -22.030 148.710 -21.790 ;
        RECT 146.410 -22.140 146.860 -22.030 ;
        RECT 148.260 -22.140 148.710 -22.030 ;
        RECT 149.920 -21.790 150.370 -21.690 ;
        RECT 150.760 -21.790 151.170 -21.360 ;
        RECT 153.920 -21.430 155.470 -21.210 ;
        RECT 155.850 -21.220 156.280 -21.160 ;
        RECT 156.660 -21.210 157.110 -21.160 ;
        RECT 157.710 -21.210 158.210 -20.820 ;
        RECT 156.660 -21.430 158.210 -21.210 ;
        RECT 167.420 -20.820 168.970 -20.600 ;
        RECT 167.420 -21.210 167.920 -20.820 ;
        RECT 168.520 -20.870 168.970 -20.820 ;
        RECT 169.350 -20.870 169.780 -20.810 ;
        RECT 170.160 -20.820 171.710 -20.600 ;
        RECT 174.460 -20.670 174.870 -20.240 ;
        RECT 175.260 -20.340 175.710 -20.240 ;
        RECT 176.920 -20.000 177.370 -19.890 ;
        RECT 178.770 -20.000 179.220 -19.890 ;
        RECT 176.920 -20.240 179.220 -20.000 ;
        RECT 176.920 -20.340 177.370 -20.240 ;
        RECT 177.760 -20.670 178.170 -20.240 ;
        RECT 178.770 -20.310 179.220 -20.240 ;
        RECT 180.170 -20.000 180.620 -19.920 ;
        RECT 181.220 -20.000 181.630 -19.560 ;
        RECT 182.020 -20.000 182.470 -19.890 ;
        RECT 180.170 -20.240 182.470 -20.000 ;
        RECT 180.170 -20.340 180.620 -20.240 ;
        RECT 182.020 -20.340 182.470 -20.240 ;
        RECT 183.660 -20.000 184.110 -19.890 ;
        RECT 184.500 -20.000 184.910 -19.560 ;
        RECT 187.680 -19.830 188.130 -19.550 ;
        RECT 191.500 -19.830 191.950 -19.550 ;
        RECT 201.180 -19.550 202.710 -19.340 ;
        RECT 203.090 -19.430 203.540 -19.340 ;
        RECT 203.920 -19.550 205.450 -19.340 ;
        RECT 185.510 -20.000 185.960 -19.920 ;
        RECT 183.660 -20.240 185.960 -20.000 ;
        RECT 183.660 -20.340 184.110 -20.240 ;
        RECT 185.510 -20.340 185.960 -20.240 ;
        RECT 186.910 -20.000 187.360 -19.890 ;
        RECT 188.760 -20.000 189.210 -19.890 ;
        RECT 186.910 -20.240 189.210 -20.000 ;
        RECT 186.910 -20.310 187.360 -20.240 ;
        RECT 170.160 -20.870 170.610 -20.820 ;
        RECT 168.520 -21.160 170.610 -20.870 ;
        RECT 168.520 -21.210 168.970 -21.160 ;
        RECT 151.770 -21.790 152.220 -21.720 ;
        RECT 149.920 -22.030 152.220 -21.790 ;
        RECT 149.920 -22.140 150.370 -22.030 ;
        RECT 151.770 -22.140 152.220 -22.030 ;
        RECT 153.170 -21.790 153.620 -21.690 ;
        RECT 155.020 -21.790 155.470 -21.690 ;
        RECT 153.170 -22.030 155.470 -21.790 ;
        RECT 153.170 -22.110 153.620 -22.030 ;
        RECT 133.680 -22.690 135.210 -22.480 ;
        RECT 135.590 -22.690 136.040 -22.600 ;
        RECT 136.420 -22.690 137.950 -22.480 ;
        RECT 147.180 -22.480 147.630 -22.200 ;
        RECT 151.000 -22.480 151.450 -22.200 ;
        RECT 154.220 -22.470 154.630 -22.030 ;
        RECT 155.020 -22.140 155.470 -22.030 ;
        RECT 156.660 -21.790 157.110 -21.690 ;
        RECT 158.510 -21.790 158.960 -21.690 ;
        RECT 156.660 -22.030 158.960 -21.790 ;
        RECT 156.660 -22.140 157.110 -22.030 ;
        RECT 157.500 -22.470 157.910 -22.030 ;
        RECT 158.510 -22.110 158.960 -22.030 ;
        RECT 159.910 -21.790 160.360 -21.720 ;
        RECT 160.960 -21.790 161.370 -21.360 ;
        RECT 161.760 -21.790 162.210 -21.690 ;
        RECT 159.910 -22.030 162.210 -21.790 ;
        RECT 159.910 -22.140 160.360 -22.030 ;
        RECT 161.760 -22.140 162.210 -22.030 ;
        RECT 163.420 -21.790 163.870 -21.690 ;
        RECT 164.260 -21.790 164.670 -21.360 ;
        RECT 167.420 -21.430 168.970 -21.210 ;
        RECT 169.350 -21.220 169.780 -21.160 ;
        RECT 170.160 -21.210 170.610 -21.160 ;
        RECT 171.210 -21.210 171.710 -20.820 ;
        RECT 170.160 -21.430 171.710 -21.210 ;
        RECT 180.920 -20.820 182.470 -20.600 ;
        RECT 180.920 -21.210 181.420 -20.820 ;
        RECT 182.020 -20.870 182.470 -20.820 ;
        RECT 182.850 -20.870 183.280 -20.810 ;
        RECT 183.660 -20.820 185.210 -20.600 ;
        RECT 187.960 -20.670 188.370 -20.240 ;
        RECT 188.760 -20.340 189.210 -20.240 ;
        RECT 190.420 -20.000 190.870 -19.890 ;
        RECT 192.270 -20.000 192.720 -19.890 ;
        RECT 190.420 -20.240 192.720 -20.000 ;
        RECT 190.420 -20.340 190.870 -20.240 ;
        RECT 191.260 -20.670 191.670 -20.240 ;
        RECT 192.270 -20.310 192.720 -20.240 ;
        RECT 193.670 -20.000 194.120 -19.920 ;
        RECT 194.720 -20.000 195.130 -19.560 ;
        RECT 195.520 -20.000 195.970 -19.890 ;
        RECT 193.670 -20.240 195.970 -20.000 ;
        RECT 193.670 -20.340 194.120 -20.240 ;
        RECT 195.520 -20.340 195.970 -20.240 ;
        RECT 197.160 -20.000 197.610 -19.890 ;
        RECT 198.000 -20.000 198.410 -19.560 ;
        RECT 201.180 -19.830 201.630 -19.550 ;
        RECT 205.000 -19.830 205.450 -19.550 ;
        RECT 214.680 -19.550 216.210 -19.340 ;
        RECT 216.590 -19.430 217.030 -19.340 ;
        RECT 199.010 -20.000 199.460 -19.920 ;
        RECT 197.160 -20.240 199.460 -20.000 ;
        RECT 197.160 -20.340 197.610 -20.240 ;
        RECT 199.010 -20.340 199.460 -20.240 ;
        RECT 200.410 -20.000 200.860 -19.890 ;
        RECT 202.260 -20.000 202.710 -19.890 ;
        RECT 200.410 -20.240 202.710 -20.000 ;
        RECT 200.410 -20.310 200.860 -20.240 ;
        RECT 183.660 -20.870 184.110 -20.820 ;
        RECT 182.020 -21.160 184.110 -20.870 ;
        RECT 182.020 -21.210 182.470 -21.160 ;
        RECT 165.270 -21.790 165.720 -21.720 ;
        RECT 163.420 -22.030 165.720 -21.790 ;
        RECT 163.420 -22.140 163.870 -22.030 ;
        RECT 165.270 -22.140 165.720 -22.030 ;
        RECT 166.670 -21.790 167.120 -21.690 ;
        RECT 168.520 -21.790 168.970 -21.690 ;
        RECT 166.670 -22.030 168.970 -21.790 ;
        RECT 166.670 -22.110 167.120 -22.030 ;
        RECT 147.180 -22.690 148.710 -22.480 ;
        RECT 149.090 -22.690 149.540 -22.600 ;
        RECT 149.920 -22.690 151.450 -22.480 ;
        RECT 160.680 -22.480 161.130 -22.200 ;
        RECT 164.500 -22.480 164.950 -22.200 ;
        RECT 167.720 -22.470 168.130 -22.030 ;
        RECT 168.520 -22.140 168.970 -22.030 ;
        RECT 170.160 -21.790 170.610 -21.690 ;
        RECT 172.010 -21.790 172.460 -21.690 ;
        RECT 170.160 -22.030 172.460 -21.790 ;
        RECT 170.160 -22.140 170.610 -22.030 ;
        RECT 171.000 -22.470 171.410 -22.030 ;
        RECT 172.010 -22.110 172.460 -22.030 ;
        RECT 173.410 -21.790 173.860 -21.720 ;
        RECT 174.460 -21.790 174.870 -21.360 ;
        RECT 175.260 -21.790 175.710 -21.690 ;
        RECT 173.410 -22.030 175.710 -21.790 ;
        RECT 173.410 -22.140 173.860 -22.030 ;
        RECT 175.260 -22.140 175.710 -22.030 ;
        RECT 176.920 -21.790 177.370 -21.690 ;
        RECT 177.760 -21.790 178.170 -21.360 ;
        RECT 180.920 -21.430 182.470 -21.210 ;
        RECT 182.850 -21.220 183.280 -21.160 ;
        RECT 183.660 -21.210 184.110 -21.160 ;
        RECT 184.710 -21.210 185.210 -20.820 ;
        RECT 183.660 -21.430 185.210 -21.210 ;
        RECT 194.420 -20.820 195.970 -20.600 ;
        RECT 194.420 -21.210 194.920 -20.820 ;
        RECT 195.520 -20.870 195.970 -20.820 ;
        RECT 196.350 -20.870 196.780 -20.810 ;
        RECT 197.160 -20.820 198.710 -20.600 ;
        RECT 201.460 -20.670 201.870 -20.240 ;
        RECT 202.260 -20.340 202.710 -20.240 ;
        RECT 203.920 -20.000 204.370 -19.890 ;
        RECT 205.770 -20.000 206.220 -19.890 ;
        RECT 203.920 -20.240 206.220 -20.000 ;
        RECT 203.920 -20.340 204.370 -20.240 ;
        RECT 204.760 -20.670 205.170 -20.240 ;
        RECT 205.770 -20.310 206.220 -20.240 ;
        RECT 207.170 -20.000 207.620 -19.920 ;
        RECT 208.220 -20.000 208.630 -19.560 ;
        RECT 209.020 -20.000 209.470 -19.890 ;
        RECT 207.170 -20.240 209.470 -20.000 ;
        RECT 207.170 -20.340 207.620 -20.240 ;
        RECT 209.020 -20.340 209.470 -20.240 ;
        RECT 210.660 -20.000 211.110 -19.890 ;
        RECT 211.500 -20.000 211.910 -19.560 ;
        RECT 214.680 -19.830 215.130 -19.550 ;
        RECT 212.510 -20.000 212.960 -19.920 ;
        RECT 210.660 -20.240 212.960 -20.000 ;
        RECT 210.660 -20.340 211.110 -20.240 ;
        RECT 212.510 -20.340 212.960 -20.240 ;
        RECT 213.910 -20.000 214.360 -19.890 ;
        RECT 215.760 -20.000 216.210 -19.890 ;
        RECT 213.910 -20.240 216.210 -20.000 ;
        RECT 213.910 -20.310 214.360 -20.240 ;
        RECT 197.160 -20.870 197.610 -20.820 ;
        RECT 195.520 -21.160 197.610 -20.870 ;
        RECT 195.520 -21.210 195.970 -21.160 ;
        RECT 178.770 -21.790 179.220 -21.720 ;
        RECT 176.920 -22.030 179.220 -21.790 ;
        RECT 176.920 -22.140 177.370 -22.030 ;
        RECT 178.770 -22.140 179.220 -22.030 ;
        RECT 180.170 -21.790 180.620 -21.690 ;
        RECT 182.020 -21.790 182.470 -21.690 ;
        RECT 180.170 -22.030 182.470 -21.790 ;
        RECT 180.170 -22.110 180.620 -22.030 ;
        RECT 160.680 -22.690 162.210 -22.480 ;
        RECT 162.590 -22.690 163.040 -22.600 ;
        RECT 163.420 -22.690 164.950 -22.480 ;
        RECT 174.180 -22.480 174.630 -22.200 ;
        RECT 178.000 -22.480 178.450 -22.200 ;
        RECT 181.220 -22.470 181.630 -22.030 ;
        RECT 182.020 -22.140 182.470 -22.030 ;
        RECT 183.660 -21.790 184.110 -21.690 ;
        RECT 185.510 -21.790 185.960 -21.690 ;
        RECT 183.660 -22.030 185.960 -21.790 ;
        RECT 183.660 -22.140 184.110 -22.030 ;
        RECT 184.500 -22.470 184.910 -22.030 ;
        RECT 185.510 -22.110 185.960 -22.030 ;
        RECT 186.910 -21.790 187.360 -21.720 ;
        RECT 187.960 -21.790 188.370 -21.360 ;
        RECT 188.760 -21.790 189.210 -21.690 ;
        RECT 186.910 -22.030 189.210 -21.790 ;
        RECT 186.910 -22.140 187.360 -22.030 ;
        RECT 188.760 -22.140 189.210 -22.030 ;
        RECT 190.420 -21.790 190.870 -21.690 ;
        RECT 191.260 -21.790 191.670 -21.360 ;
        RECT 194.420 -21.430 195.970 -21.210 ;
        RECT 196.350 -21.220 196.780 -21.160 ;
        RECT 197.160 -21.210 197.610 -21.160 ;
        RECT 198.210 -21.210 198.710 -20.820 ;
        RECT 197.160 -21.430 198.710 -21.210 ;
        RECT 207.920 -20.820 209.470 -20.600 ;
        RECT 207.920 -21.210 208.420 -20.820 ;
        RECT 209.020 -20.870 209.470 -20.820 ;
        RECT 209.850 -20.870 210.280 -20.810 ;
        RECT 210.660 -20.820 212.210 -20.600 ;
        RECT 214.960 -20.670 215.370 -20.240 ;
        RECT 215.760 -20.340 216.210 -20.240 ;
        RECT 210.660 -20.870 211.110 -20.820 ;
        RECT 209.020 -21.160 211.110 -20.870 ;
        RECT 209.020 -21.210 209.470 -21.160 ;
        RECT 192.270 -21.790 192.720 -21.720 ;
        RECT 190.420 -22.030 192.720 -21.790 ;
        RECT 190.420 -22.140 190.870 -22.030 ;
        RECT 192.270 -22.140 192.720 -22.030 ;
        RECT 193.670 -21.790 194.120 -21.690 ;
        RECT 195.520 -21.790 195.970 -21.690 ;
        RECT 193.670 -22.030 195.970 -21.790 ;
        RECT 193.670 -22.110 194.120 -22.030 ;
        RECT 174.180 -22.690 175.710 -22.480 ;
        RECT 176.090 -22.690 176.540 -22.600 ;
        RECT 176.920 -22.690 178.450 -22.480 ;
        RECT 187.680 -22.480 188.130 -22.200 ;
        RECT 191.500 -22.480 191.950 -22.200 ;
        RECT 194.720 -22.470 195.130 -22.030 ;
        RECT 195.520 -22.140 195.970 -22.030 ;
        RECT 197.160 -21.790 197.610 -21.690 ;
        RECT 199.010 -21.790 199.460 -21.690 ;
        RECT 197.160 -22.030 199.460 -21.790 ;
        RECT 197.160 -22.140 197.610 -22.030 ;
        RECT 198.000 -22.470 198.410 -22.030 ;
        RECT 199.010 -22.110 199.460 -22.030 ;
        RECT 200.410 -21.790 200.860 -21.720 ;
        RECT 201.460 -21.790 201.870 -21.360 ;
        RECT 202.260 -21.790 202.710 -21.690 ;
        RECT 200.410 -22.030 202.710 -21.790 ;
        RECT 200.410 -22.140 200.860 -22.030 ;
        RECT 202.260 -22.140 202.710 -22.030 ;
        RECT 203.920 -21.790 204.370 -21.690 ;
        RECT 204.760 -21.790 205.170 -21.360 ;
        RECT 207.920 -21.430 209.470 -21.210 ;
        RECT 209.850 -21.220 210.280 -21.160 ;
        RECT 210.660 -21.210 211.110 -21.160 ;
        RECT 211.710 -21.210 212.210 -20.820 ;
        RECT 210.660 -21.430 212.210 -21.210 ;
        RECT 205.770 -21.790 206.220 -21.720 ;
        RECT 203.920 -22.030 206.220 -21.790 ;
        RECT 203.920 -22.140 204.370 -22.030 ;
        RECT 205.770 -22.140 206.220 -22.030 ;
        RECT 207.170 -21.790 207.620 -21.690 ;
        RECT 209.020 -21.790 209.470 -21.690 ;
        RECT 207.170 -22.030 209.470 -21.790 ;
        RECT 207.170 -22.110 207.620 -22.030 ;
        RECT 187.680 -22.690 189.210 -22.480 ;
        RECT 189.590 -22.690 190.040 -22.600 ;
        RECT 190.420 -22.690 191.950 -22.480 ;
        RECT 201.180 -22.480 201.630 -22.200 ;
        RECT 205.000 -22.480 205.450 -22.200 ;
        RECT 208.220 -22.470 208.630 -22.030 ;
        RECT 209.020 -22.140 209.470 -22.030 ;
        RECT 210.660 -21.790 211.110 -21.690 ;
        RECT 212.510 -21.790 212.960 -21.690 ;
        RECT 210.660 -22.030 212.960 -21.790 ;
        RECT 210.660 -22.140 211.110 -22.030 ;
        RECT 211.500 -22.470 211.910 -22.030 ;
        RECT 212.510 -22.110 212.960 -22.030 ;
        RECT 213.910 -21.790 214.360 -21.720 ;
        RECT 214.960 -21.790 215.370 -21.360 ;
        RECT 215.760 -21.790 216.210 -21.690 ;
        RECT 213.910 -22.030 216.210 -21.790 ;
        RECT 213.910 -22.140 214.360 -22.030 ;
        RECT 215.760 -22.140 216.210 -22.030 ;
        RECT 201.180 -22.690 202.710 -22.480 ;
        RECT 203.090 -22.690 203.540 -22.600 ;
        RECT 203.920 -22.690 205.450 -22.480 ;
        RECT 214.680 -22.480 215.130 -22.200 ;
        RECT 214.680 -22.690 216.210 -22.480 ;
        RECT 216.590 -22.690 217.030 -22.600 ;
        RECT 13.260 -22.950 15.370 -22.690 ;
        RECT 26.760 -22.950 28.870 -22.690 ;
        RECT 40.260 -22.950 42.370 -22.690 ;
        RECT 53.760 -22.950 55.870 -22.690 ;
        RECT 67.260 -22.950 69.370 -22.690 ;
        RECT 80.760 -22.950 82.870 -22.690 ;
        RECT 94.260 -22.950 96.370 -22.690 ;
        RECT 107.760 -22.950 109.870 -22.690 ;
        RECT 121.260 -22.950 123.370 -22.690 ;
        RECT 134.760 -22.950 136.870 -22.690 ;
        RECT 148.260 -22.950 150.370 -22.690 ;
        RECT 161.760 -22.950 163.870 -22.690 ;
        RECT 175.260 -22.950 177.370 -22.690 ;
        RECT 188.760 -22.950 190.870 -22.690 ;
        RECT 202.260 -22.950 204.370 -22.690 ;
        RECT 215.760 -22.750 217.030 -22.690 ;
        RECT 215.760 -22.940 217.240 -22.750 ;
        RECT 215.760 -22.950 217.030 -22.940 ;
        RECT 12.180 -23.160 13.710 -22.950 ;
        RECT 14.090 -23.040 14.540 -22.950 ;
        RECT 14.920 -23.160 16.450 -22.950 ;
        RECT 1.420 -23.610 1.870 -23.500 ;
        RECT 3.270 -23.610 3.720 -23.500 ;
        RECT 1.420 -23.850 3.720 -23.610 ;
        RECT 1.420 -23.950 1.870 -23.850 ;
        RECT 2.260 -24.280 2.670 -23.850 ;
        RECT 3.270 -23.920 3.720 -23.850 ;
        RECT 4.670 -23.610 5.120 -23.530 ;
        RECT 5.720 -23.610 6.130 -23.170 ;
        RECT 6.520 -23.610 6.970 -23.500 ;
        RECT 4.670 -23.850 6.970 -23.610 ;
        RECT 4.670 -23.950 5.120 -23.850 ;
        RECT 6.520 -23.950 6.970 -23.850 ;
        RECT 8.160 -23.610 8.610 -23.500 ;
        RECT 9.000 -23.610 9.410 -23.170 ;
        RECT 12.180 -23.440 12.630 -23.160 ;
        RECT 16.000 -23.440 16.450 -23.160 ;
        RECT 25.680 -23.160 27.210 -22.950 ;
        RECT 27.590 -23.040 28.040 -22.950 ;
        RECT 28.420 -23.160 29.950 -22.950 ;
        RECT 10.010 -23.610 10.460 -23.530 ;
        RECT 8.160 -23.850 10.460 -23.610 ;
        RECT 8.160 -23.950 8.610 -23.850 ;
        RECT 10.010 -23.950 10.460 -23.850 ;
        RECT 11.410 -23.610 11.860 -23.500 ;
        RECT 13.260 -23.610 13.710 -23.500 ;
        RECT 11.410 -23.850 13.710 -23.610 ;
        RECT 11.410 -23.920 11.860 -23.850 ;
        RECT 5.420 -24.430 6.970 -24.210 ;
        RECT 5.420 -24.820 5.920 -24.430 ;
        RECT 6.520 -24.480 6.970 -24.430 ;
        RECT 7.350 -24.480 7.780 -24.420 ;
        RECT 8.160 -24.430 9.710 -24.210 ;
        RECT 12.460 -24.280 12.870 -23.850 ;
        RECT 13.260 -23.950 13.710 -23.850 ;
        RECT 14.920 -23.610 15.370 -23.500 ;
        RECT 16.770 -23.610 17.220 -23.500 ;
        RECT 14.920 -23.850 17.220 -23.610 ;
        RECT 14.920 -23.950 15.370 -23.850 ;
        RECT 15.760 -24.280 16.170 -23.850 ;
        RECT 16.770 -23.920 17.220 -23.850 ;
        RECT 18.170 -23.610 18.620 -23.530 ;
        RECT 19.220 -23.610 19.630 -23.170 ;
        RECT 20.020 -23.610 20.470 -23.500 ;
        RECT 18.170 -23.850 20.470 -23.610 ;
        RECT 18.170 -23.950 18.620 -23.850 ;
        RECT 20.020 -23.950 20.470 -23.850 ;
        RECT 21.660 -23.610 22.110 -23.500 ;
        RECT 22.500 -23.610 22.910 -23.170 ;
        RECT 25.680 -23.440 26.130 -23.160 ;
        RECT 29.500 -23.440 29.950 -23.160 ;
        RECT 39.180 -23.160 40.710 -22.950 ;
        RECT 41.090 -23.040 41.540 -22.950 ;
        RECT 41.920 -23.160 43.450 -22.950 ;
        RECT 23.510 -23.610 23.960 -23.530 ;
        RECT 21.660 -23.850 23.960 -23.610 ;
        RECT 21.660 -23.950 22.110 -23.850 ;
        RECT 23.510 -23.950 23.960 -23.850 ;
        RECT 24.910 -23.610 25.360 -23.500 ;
        RECT 26.760 -23.610 27.210 -23.500 ;
        RECT 24.910 -23.850 27.210 -23.610 ;
        RECT 24.910 -23.920 25.360 -23.850 ;
        RECT 8.160 -24.480 8.610 -24.430 ;
        RECT 6.520 -24.770 8.610 -24.480 ;
        RECT 6.520 -24.820 6.970 -24.770 ;
        RECT 1.420 -25.400 1.870 -25.300 ;
        RECT 2.260 -25.400 2.670 -24.970 ;
        RECT 5.420 -25.040 6.970 -24.820 ;
        RECT 7.350 -24.830 7.780 -24.770 ;
        RECT 8.160 -24.820 8.610 -24.770 ;
        RECT 9.210 -24.820 9.710 -24.430 ;
        RECT 8.160 -25.040 9.710 -24.820 ;
        RECT 18.920 -24.430 20.470 -24.210 ;
        RECT 18.920 -24.820 19.420 -24.430 ;
        RECT 20.020 -24.480 20.470 -24.430 ;
        RECT 20.850 -24.480 21.280 -24.420 ;
        RECT 21.660 -24.430 23.210 -24.210 ;
        RECT 25.960 -24.280 26.370 -23.850 ;
        RECT 26.760 -23.950 27.210 -23.850 ;
        RECT 28.420 -23.610 28.870 -23.500 ;
        RECT 30.270 -23.610 30.720 -23.500 ;
        RECT 28.420 -23.850 30.720 -23.610 ;
        RECT 28.420 -23.950 28.870 -23.850 ;
        RECT 29.260 -24.280 29.670 -23.850 ;
        RECT 30.270 -23.920 30.720 -23.850 ;
        RECT 31.670 -23.610 32.120 -23.530 ;
        RECT 32.720 -23.610 33.130 -23.170 ;
        RECT 33.520 -23.610 33.970 -23.500 ;
        RECT 31.670 -23.850 33.970 -23.610 ;
        RECT 31.670 -23.950 32.120 -23.850 ;
        RECT 33.520 -23.950 33.970 -23.850 ;
        RECT 35.160 -23.610 35.610 -23.500 ;
        RECT 36.000 -23.610 36.410 -23.170 ;
        RECT 39.180 -23.440 39.630 -23.160 ;
        RECT 43.000 -23.440 43.450 -23.160 ;
        RECT 52.680 -23.160 54.210 -22.950 ;
        RECT 54.590 -23.040 55.040 -22.950 ;
        RECT 55.420 -23.160 56.950 -22.950 ;
        RECT 37.010 -23.610 37.460 -23.530 ;
        RECT 35.160 -23.850 37.460 -23.610 ;
        RECT 35.160 -23.950 35.610 -23.850 ;
        RECT 37.010 -23.950 37.460 -23.850 ;
        RECT 38.410 -23.610 38.860 -23.500 ;
        RECT 40.260 -23.610 40.710 -23.500 ;
        RECT 38.410 -23.850 40.710 -23.610 ;
        RECT 38.410 -23.920 38.860 -23.850 ;
        RECT 21.660 -24.480 22.110 -24.430 ;
        RECT 20.020 -24.770 22.110 -24.480 ;
        RECT 20.020 -24.820 20.470 -24.770 ;
        RECT 3.270 -25.400 3.720 -25.330 ;
        RECT 1.420 -25.640 3.720 -25.400 ;
        RECT 1.420 -25.750 1.870 -25.640 ;
        RECT 3.270 -25.750 3.720 -25.640 ;
        RECT 4.670 -25.400 5.120 -25.300 ;
        RECT 6.520 -25.400 6.970 -25.300 ;
        RECT 4.670 -25.640 6.970 -25.400 ;
        RECT 4.670 -25.720 5.120 -25.640 ;
        RECT 5.720 -26.080 6.130 -25.640 ;
        RECT 6.520 -25.750 6.970 -25.640 ;
        RECT 8.160 -25.400 8.610 -25.300 ;
        RECT 10.010 -25.400 10.460 -25.300 ;
        RECT 8.160 -25.640 10.460 -25.400 ;
        RECT 8.160 -25.750 8.610 -25.640 ;
        RECT 9.000 -26.080 9.410 -25.640 ;
        RECT 10.010 -25.720 10.460 -25.640 ;
        RECT 11.410 -25.400 11.860 -25.330 ;
        RECT 12.460 -25.400 12.870 -24.970 ;
        RECT 13.260 -25.400 13.710 -25.300 ;
        RECT 11.410 -25.640 13.710 -25.400 ;
        RECT 11.410 -25.750 11.860 -25.640 ;
        RECT 13.260 -25.750 13.710 -25.640 ;
        RECT 14.920 -25.400 15.370 -25.300 ;
        RECT 15.760 -25.400 16.170 -24.970 ;
        RECT 18.920 -25.040 20.470 -24.820 ;
        RECT 20.850 -24.830 21.280 -24.770 ;
        RECT 21.660 -24.820 22.110 -24.770 ;
        RECT 22.710 -24.820 23.210 -24.430 ;
        RECT 21.660 -25.040 23.210 -24.820 ;
        RECT 32.420 -24.430 33.970 -24.210 ;
        RECT 32.420 -24.820 32.920 -24.430 ;
        RECT 33.520 -24.480 33.970 -24.430 ;
        RECT 34.350 -24.480 34.780 -24.420 ;
        RECT 35.160 -24.430 36.710 -24.210 ;
        RECT 39.460 -24.280 39.870 -23.850 ;
        RECT 40.260 -23.950 40.710 -23.850 ;
        RECT 41.920 -23.610 42.370 -23.500 ;
        RECT 43.770 -23.610 44.220 -23.500 ;
        RECT 41.920 -23.850 44.220 -23.610 ;
        RECT 41.920 -23.950 42.370 -23.850 ;
        RECT 42.760 -24.280 43.170 -23.850 ;
        RECT 43.770 -23.920 44.220 -23.850 ;
        RECT 45.170 -23.610 45.620 -23.530 ;
        RECT 46.220 -23.610 46.630 -23.170 ;
        RECT 47.020 -23.610 47.470 -23.500 ;
        RECT 45.170 -23.850 47.470 -23.610 ;
        RECT 45.170 -23.950 45.620 -23.850 ;
        RECT 47.020 -23.950 47.470 -23.850 ;
        RECT 48.660 -23.610 49.110 -23.500 ;
        RECT 49.500 -23.610 49.910 -23.170 ;
        RECT 52.680 -23.440 53.130 -23.160 ;
        RECT 56.500 -23.440 56.950 -23.160 ;
        RECT 66.180 -23.160 67.710 -22.950 ;
        RECT 68.090 -23.040 68.540 -22.950 ;
        RECT 68.920 -23.160 70.450 -22.950 ;
        RECT 50.510 -23.610 50.960 -23.530 ;
        RECT 48.660 -23.850 50.960 -23.610 ;
        RECT 48.660 -23.950 49.110 -23.850 ;
        RECT 50.510 -23.950 50.960 -23.850 ;
        RECT 51.910 -23.610 52.360 -23.500 ;
        RECT 53.760 -23.610 54.210 -23.500 ;
        RECT 51.910 -23.850 54.210 -23.610 ;
        RECT 51.910 -23.920 52.360 -23.850 ;
        RECT 35.160 -24.480 35.610 -24.430 ;
        RECT 33.520 -24.770 35.610 -24.480 ;
        RECT 33.520 -24.820 33.970 -24.770 ;
        RECT 16.770 -25.400 17.220 -25.330 ;
        RECT 14.920 -25.640 17.220 -25.400 ;
        RECT 14.920 -25.750 15.370 -25.640 ;
        RECT 16.770 -25.750 17.220 -25.640 ;
        RECT 18.170 -25.400 18.620 -25.300 ;
        RECT 20.020 -25.400 20.470 -25.300 ;
        RECT 18.170 -25.640 20.470 -25.400 ;
        RECT 18.170 -25.720 18.620 -25.640 ;
        RECT 12.180 -26.090 12.630 -25.810 ;
        RECT 16.000 -26.090 16.450 -25.810 ;
        RECT 19.220 -26.080 19.630 -25.640 ;
        RECT 20.020 -25.750 20.470 -25.640 ;
        RECT 21.660 -25.400 22.110 -25.300 ;
        RECT 23.510 -25.400 23.960 -25.300 ;
        RECT 21.660 -25.640 23.960 -25.400 ;
        RECT 21.660 -25.750 22.110 -25.640 ;
        RECT 22.500 -26.080 22.910 -25.640 ;
        RECT 23.510 -25.720 23.960 -25.640 ;
        RECT 24.910 -25.400 25.360 -25.330 ;
        RECT 25.960 -25.400 26.370 -24.970 ;
        RECT 26.760 -25.400 27.210 -25.300 ;
        RECT 24.910 -25.640 27.210 -25.400 ;
        RECT 24.910 -25.750 25.360 -25.640 ;
        RECT 26.760 -25.750 27.210 -25.640 ;
        RECT 28.420 -25.400 28.870 -25.300 ;
        RECT 29.260 -25.400 29.670 -24.970 ;
        RECT 32.420 -25.040 33.970 -24.820 ;
        RECT 34.350 -24.830 34.780 -24.770 ;
        RECT 35.160 -24.820 35.610 -24.770 ;
        RECT 36.210 -24.820 36.710 -24.430 ;
        RECT 35.160 -25.040 36.710 -24.820 ;
        RECT 45.920 -24.430 47.470 -24.210 ;
        RECT 45.920 -24.820 46.420 -24.430 ;
        RECT 47.020 -24.480 47.470 -24.430 ;
        RECT 47.850 -24.480 48.280 -24.420 ;
        RECT 48.660 -24.430 50.210 -24.210 ;
        RECT 52.960 -24.280 53.370 -23.850 ;
        RECT 53.760 -23.950 54.210 -23.850 ;
        RECT 55.420 -23.610 55.870 -23.500 ;
        RECT 57.270 -23.610 57.720 -23.500 ;
        RECT 55.420 -23.850 57.720 -23.610 ;
        RECT 55.420 -23.950 55.870 -23.850 ;
        RECT 56.260 -24.280 56.670 -23.850 ;
        RECT 57.270 -23.920 57.720 -23.850 ;
        RECT 58.670 -23.610 59.120 -23.530 ;
        RECT 59.720 -23.610 60.130 -23.170 ;
        RECT 60.520 -23.610 60.970 -23.500 ;
        RECT 58.670 -23.850 60.970 -23.610 ;
        RECT 58.670 -23.950 59.120 -23.850 ;
        RECT 60.520 -23.950 60.970 -23.850 ;
        RECT 62.160 -23.610 62.610 -23.500 ;
        RECT 63.000 -23.610 63.410 -23.170 ;
        RECT 66.180 -23.440 66.630 -23.160 ;
        RECT 70.000 -23.440 70.450 -23.160 ;
        RECT 79.680 -23.160 81.210 -22.950 ;
        RECT 81.590 -23.040 82.040 -22.950 ;
        RECT 82.420 -23.160 83.950 -22.950 ;
        RECT 64.010 -23.610 64.460 -23.530 ;
        RECT 62.160 -23.850 64.460 -23.610 ;
        RECT 62.160 -23.950 62.610 -23.850 ;
        RECT 64.010 -23.950 64.460 -23.850 ;
        RECT 65.410 -23.610 65.860 -23.500 ;
        RECT 67.260 -23.610 67.710 -23.500 ;
        RECT 65.410 -23.850 67.710 -23.610 ;
        RECT 65.410 -23.920 65.860 -23.850 ;
        RECT 48.660 -24.480 49.110 -24.430 ;
        RECT 47.020 -24.770 49.110 -24.480 ;
        RECT 47.020 -24.820 47.470 -24.770 ;
        RECT 30.270 -25.400 30.720 -25.330 ;
        RECT 28.420 -25.640 30.720 -25.400 ;
        RECT 28.420 -25.750 28.870 -25.640 ;
        RECT 30.270 -25.750 30.720 -25.640 ;
        RECT 31.670 -25.400 32.120 -25.300 ;
        RECT 33.520 -25.400 33.970 -25.300 ;
        RECT 31.670 -25.640 33.970 -25.400 ;
        RECT 31.670 -25.720 32.120 -25.640 ;
        RECT 12.180 -26.300 13.710 -26.090 ;
        RECT 14.090 -26.300 14.540 -26.210 ;
        RECT 14.920 -26.300 16.450 -26.090 ;
        RECT 25.680 -26.090 26.130 -25.810 ;
        RECT 29.500 -26.090 29.950 -25.810 ;
        RECT 32.720 -26.080 33.130 -25.640 ;
        RECT 33.520 -25.750 33.970 -25.640 ;
        RECT 35.160 -25.400 35.610 -25.300 ;
        RECT 37.010 -25.400 37.460 -25.300 ;
        RECT 35.160 -25.640 37.460 -25.400 ;
        RECT 35.160 -25.750 35.610 -25.640 ;
        RECT 36.000 -26.080 36.410 -25.640 ;
        RECT 37.010 -25.720 37.460 -25.640 ;
        RECT 38.410 -25.400 38.860 -25.330 ;
        RECT 39.460 -25.400 39.870 -24.970 ;
        RECT 40.260 -25.400 40.710 -25.300 ;
        RECT 38.410 -25.640 40.710 -25.400 ;
        RECT 38.410 -25.750 38.860 -25.640 ;
        RECT 40.260 -25.750 40.710 -25.640 ;
        RECT 41.920 -25.400 42.370 -25.300 ;
        RECT 42.760 -25.400 43.170 -24.970 ;
        RECT 45.920 -25.040 47.470 -24.820 ;
        RECT 47.850 -24.830 48.280 -24.770 ;
        RECT 48.660 -24.820 49.110 -24.770 ;
        RECT 49.710 -24.820 50.210 -24.430 ;
        RECT 48.660 -25.040 50.210 -24.820 ;
        RECT 59.420 -24.430 60.970 -24.210 ;
        RECT 59.420 -24.820 59.920 -24.430 ;
        RECT 60.520 -24.480 60.970 -24.430 ;
        RECT 61.350 -24.480 61.780 -24.420 ;
        RECT 62.160 -24.430 63.710 -24.210 ;
        RECT 66.460 -24.280 66.870 -23.850 ;
        RECT 67.260 -23.950 67.710 -23.850 ;
        RECT 68.920 -23.610 69.370 -23.500 ;
        RECT 70.770 -23.610 71.220 -23.500 ;
        RECT 68.920 -23.850 71.220 -23.610 ;
        RECT 68.920 -23.950 69.370 -23.850 ;
        RECT 69.760 -24.280 70.170 -23.850 ;
        RECT 70.770 -23.920 71.220 -23.850 ;
        RECT 72.170 -23.610 72.620 -23.530 ;
        RECT 73.220 -23.610 73.630 -23.170 ;
        RECT 74.020 -23.610 74.470 -23.500 ;
        RECT 72.170 -23.850 74.470 -23.610 ;
        RECT 72.170 -23.950 72.620 -23.850 ;
        RECT 74.020 -23.950 74.470 -23.850 ;
        RECT 75.660 -23.610 76.110 -23.500 ;
        RECT 76.500 -23.610 76.910 -23.170 ;
        RECT 79.680 -23.440 80.130 -23.160 ;
        RECT 83.500 -23.440 83.950 -23.160 ;
        RECT 93.180 -23.160 94.710 -22.950 ;
        RECT 95.090 -23.040 95.540 -22.950 ;
        RECT 95.920 -23.160 97.450 -22.950 ;
        RECT 77.510 -23.610 77.960 -23.530 ;
        RECT 75.660 -23.850 77.960 -23.610 ;
        RECT 75.660 -23.950 76.110 -23.850 ;
        RECT 77.510 -23.950 77.960 -23.850 ;
        RECT 78.910 -23.610 79.360 -23.500 ;
        RECT 80.760 -23.610 81.210 -23.500 ;
        RECT 78.910 -23.850 81.210 -23.610 ;
        RECT 78.910 -23.920 79.360 -23.850 ;
        RECT 62.160 -24.480 62.610 -24.430 ;
        RECT 60.520 -24.770 62.610 -24.480 ;
        RECT 60.520 -24.820 60.970 -24.770 ;
        RECT 43.770 -25.400 44.220 -25.330 ;
        RECT 41.920 -25.640 44.220 -25.400 ;
        RECT 41.920 -25.750 42.370 -25.640 ;
        RECT 43.770 -25.750 44.220 -25.640 ;
        RECT 45.170 -25.400 45.620 -25.300 ;
        RECT 47.020 -25.400 47.470 -25.300 ;
        RECT 45.170 -25.640 47.470 -25.400 ;
        RECT 45.170 -25.720 45.620 -25.640 ;
        RECT 25.680 -26.300 27.210 -26.090 ;
        RECT 27.590 -26.300 28.040 -26.210 ;
        RECT 28.420 -26.300 29.950 -26.090 ;
        RECT 39.180 -26.090 39.630 -25.810 ;
        RECT 43.000 -26.090 43.450 -25.810 ;
        RECT 46.220 -26.080 46.630 -25.640 ;
        RECT 47.020 -25.750 47.470 -25.640 ;
        RECT 48.660 -25.400 49.110 -25.300 ;
        RECT 50.510 -25.400 50.960 -25.300 ;
        RECT 48.660 -25.640 50.960 -25.400 ;
        RECT 48.660 -25.750 49.110 -25.640 ;
        RECT 49.500 -26.080 49.910 -25.640 ;
        RECT 50.510 -25.720 50.960 -25.640 ;
        RECT 51.910 -25.400 52.360 -25.330 ;
        RECT 52.960 -25.400 53.370 -24.970 ;
        RECT 53.760 -25.400 54.210 -25.300 ;
        RECT 51.910 -25.640 54.210 -25.400 ;
        RECT 51.910 -25.750 52.360 -25.640 ;
        RECT 53.760 -25.750 54.210 -25.640 ;
        RECT 55.420 -25.400 55.870 -25.300 ;
        RECT 56.260 -25.400 56.670 -24.970 ;
        RECT 59.420 -25.040 60.970 -24.820 ;
        RECT 61.350 -24.830 61.780 -24.770 ;
        RECT 62.160 -24.820 62.610 -24.770 ;
        RECT 63.210 -24.820 63.710 -24.430 ;
        RECT 62.160 -25.040 63.710 -24.820 ;
        RECT 72.920 -24.430 74.470 -24.210 ;
        RECT 72.920 -24.820 73.420 -24.430 ;
        RECT 74.020 -24.480 74.470 -24.430 ;
        RECT 74.850 -24.480 75.280 -24.420 ;
        RECT 75.660 -24.430 77.210 -24.210 ;
        RECT 79.960 -24.280 80.370 -23.850 ;
        RECT 80.760 -23.950 81.210 -23.850 ;
        RECT 82.420 -23.610 82.870 -23.500 ;
        RECT 84.270 -23.610 84.720 -23.500 ;
        RECT 82.420 -23.850 84.720 -23.610 ;
        RECT 82.420 -23.950 82.870 -23.850 ;
        RECT 83.260 -24.280 83.670 -23.850 ;
        RECT 84.270 -23.920 84.720 -23.850 ;
        RECT 85.670 -23.610 86.120 -23.530 ;
        RECT 86.720 -23.610 87.130 -23.170 ;
        RECT 87.520 -23.610 87.970 -23.500 ;
        RECT 85.670 -23.850 87.970 -23.610 ;
        RECT 85.670 -23.950 86.120 -23.850 ;
        RECT 87.520 -23.950 87.970 -23.850 ;
        RECT 89.160 -23.610 89.610 -23.500 ;
        RECT 90.000 -23.610 90.410 -23.170 ;
        RECT 93.180 -23.440 93.630 -23.160 ;
        RECT 97.000 -23.440 97.450 -23.160 ;
        RECT 106.680 -23.160 108.210 -22.950 ;
        RECT 108.590 -23.040 109.040 -22.950 ;
        RECT 109.420 -23.160 110.950 -22.950 ;
        RECT 91.010 -23.610 91.460 -23.530 ;
        RECT 89.160 -23.850 91.460 -23.610 ;
        RECT 89.160 -23.950 89.610 -23.850 ;
        RECT 91.010 -23.950 91.460 -23.850 ;
        RECT 92.410 -23.610 92.860 -23.500 ;
        RECT 94.260 -23.610 94.710 -23.500 ;
        RECT 92.410 -23.850 94.710 -23.610 ;
        RECT 92.410 -23.920 92.860 -23.850 ;
        RECT 75.660 -24.480 76.110 -24.430 ;
        RECT 74.020 -24.770 76.110 -24.480 ;
        RECT 74.020 -24.820 74.470 -24.770 ;
        RECT 57.270 -25.400 57.720 -25.330 ;
        RECT 55.420 -25.640 57.720 -25.400 ;
        RECT 55.420 -25.750 55.870 -25.640 ;
        RECT 57.270 -25.750 57.720 -25.640 ;
        RECT 58.670 -25.400 59.120 -25.300 ;
        RECT 60.520 -25.400 60.970 -25.300 ;
        RECT 58.670 -25.640 60.970 -25.400 ;
        RECT 58.670 -25.720 59.120 -25.640 ;
        RECT 39.180 -26.300 40.710 -26.090 ;
        RECT 41.090 -26.300 41.540 -26.210 ;
        RECT 41.920 -26.300 43.450 -26.090 ;
        RECT 52.680 -26.090 53.130 -25.810 ;
        RECT 56.500 -26.090 56.950 -25.810 ;
        RECT 59.720 -26.080 60.130 -25.640 ;
        RECT 60.520 -25.750 60.970 -25.640 ;
        RECT 62.160 -25.400 62.610 -25.300 ;
        RECT 64.010 -25.400 64.460 -25.300 ;
        RECT 62.160 -25.640 64.460 -25.400 ;
        RECT 62.160 -25.750 62.610 -25.640 ;
        RECT 63.000 -26.080 63.410 -25.640 ;
        RECT 64.010 -25.720 64.460 -25.640 ;
        RECT 65.410 -25.400 65.860 -25.330 ;
        RECT 66.460 -25.400 66.870 -24.970 ;
        RECT 67.260 -25.400 67.710 -25.300 ;
        RECT 65.410 -25.640 67.710 -25.400 ;
        RECT 65.410 -25.750 65.860 -25.640 ;
        RECT 67.260 -25.750 67.710 -25.640 ;
        RECT 68.920 -25.400 69.370 -25.300 ;
        RECT 69.760 -25.400 70.170 -24.970 ;
        RECT 72.920 -25.040 74.470 -24.820 ;
        RECT 74.850 -24.830 75.280 -24.770 ;
        RECT 75.660 -24.820 76.110 -24.770 ;
        RECT 76.710 -24.820 77.210 -24.430 ;
        RECT 75.660 -25.040 77.210 -24.820 ;
        RECT 86.420 -24.430 87.970 -24.210 ;
        RECT 86.420 -24.820 86.920 -24.430 ;
        RECT 87.520 -24.480 87.970 -24.430 ;
        RECT 88.350 -24.480 88.780 -24.420 ;
        RECT 89.160 -24.430 90.710 -24.210 ;
        RECT 93.460 -24.280 93.870 -23.850 ;
        RECT 94.260 -23.950 94.710 -23.850 ;
        RECT 95.920 -23.610 96.370 -23.500 ;
        RECT 97.770 -23.610 98.220 -23.500 ;
        RECT 95.920 -23.850 98.220 -23.610 ;
        RECT 95.920 -23.950 96.370 -23.850 ;
        RECT 96.760 -24.280 97.170 -23.850 ;
        RECT 97.770 -23.920 98.220 -23.850 ;
        RECT 99.170 -23.610 99.620 -23.530 ;
        RECT 100.220 -23.610 100.630 -23.170 ;
        RECT 101.020 -23.610 101.470 -23.500 ;
        RECT 99.170 -23.850 101.470 -23.610 ;
        RECT 99.170 -23.950 99.620 -23.850 ;
        RECT 101.020 -23.950 101.470 -23.850 ;
        RECT 102.660 -23.610 103.110 -23.500 ;
        RECT 103.500 -23.610 103.910 -23.170 ;
        RECT 106.680 -23.440 107.130 -23.160 ;
        RECT 110.500 -23.440 110.950 -23.160 ;
        RECT 120.180 -23.160 121.710 -22.950 ;
        RECT 122.090 -23.040 122.540 -22.950 ;
        RECT 122.920 -23.160 124.450 -22.950 ;
        RECT 104.510 -23.610 104.960 -23.530 ;
        RECT 102.660 -23.850 104.960 -23.610 ;
        RECT 102.660 -23.950 103.110 -23.850 ;
        RECT 104.510 -23.950 104.960 -23.850 ;
        RECT 105.910 -23.610 106.360 -23.500 ;
        RECT 107.760 -23.610 108.210 -23.500 ;
        RECT 105.910 -23.850 108.210 -23.610 ;
        RECT 105.910 -23.920 106.360 -23.850 ;
        RECT 89.160 -24.480 89.610 -24.430 ;
        RECT 87.520 -24.770 89.610 -24.480 ;
        RECT 87.520 -24.820 87.970 -24.770 ;
        RECT 70.770 -25.400 71.220 -25.330 ;
        RECT 68.920 -25.640 71.220 -25.400 ;
        RECT 68.920 -25.750 69.370 -25.640 ;
        RECT 70.770 -25.750 71.220 -25.640 ;
        RECT 72.170 -25.400 72.620 -25.300 ;
        RECT 74.020 -25.400 74.470 -25.300 ;
        RECT 72.170 -25.640 74.470 -25.400 ;
        RECT 72.170 -25.720 72.620 -25.640 ;
        RECT 52.680 -26.250 54.210 -26.090 ;
        RECT 54.590 -26.250 55.040 -26.210 ;
        RECT 55.420 -26.250 56.950 -26.090 ;
        RECT 52.680 -26.300 56.950 -26.250 ;
        RECT 66.180 -26.090 66.630 -25.810 ;
        RECT 70.000 -26.090 70.450 -25.810 ;
        RECT 73.220 -26.080 73.630 -25.640 ;
        RECT 74.020 -25.750 74.470 -25.640 ;
        RECT 75.660 -25.400 76.110 -25.300 ;
        RECT 77.510 -25.400 77.960 -25.300 ;
        RECT 75.660 -25.640 77.960 -25.400 ;
        RECT 75.660 -25.750 76.110 -25.640 ;
        RECT 76.500 -26.080 76.910 -25.640 ;
        RECT 77.510 -25.720 77.960 -25.640 ;
        RECT 78.910 -25.400 79.360 -25.330 ;
        RECT 79.960 -25.400 80.370 -24.970 ;
        RECT 80.760 -25.400 81.210 -25.300 ;
        RECT 78.910 -25.640 81.210 -25.400 ;
        RECT 78.910 -25.750 79.360 -25.640 ;
        RECT 80.760 -25.750 81.210 -25.640 ;
        RECT 82.420 -25.400 82.870 -25.300 ;
        RECT 83.260 -25.400 83.670 -24.970 ;
        RECT 86.420 -25.040 87.970 -24.820 ;
        RECT 88.350 -24.830 88.780 -24.770 ;
        RECT 89.160 -24.820 89.610 -24.770 ;
        RECT 90.210 -24.820 90.710 -24.430 ;
        RECT 89.160 -25.040 90.710 -24.820 ;
        RECT 99.920 -24.430 101.470 -24.210 ;
        RECT 99.920 -24.820 100.420 -24.430 ;
        RECT 101.020 -24.480 101.470 -24.430 ;
        RECT 101.850 -24.480 102.280 -24.420 ;
        RECT 102.660 -24.430 104.210 -24.210 ;
        RECT 106.960 -24.280 107.370 -23.850 ;
        RECT 107.760 -23.950 108.210 -23.850 ;
        RECT 109.420 -23.610 109.870 -23.500 ;
        RECT 111.270 -23.610 111.720 -23.500 ;
        RECT 109.420 -23.850 111.720 -23.610 ;
        RECT 109.420 -23.950 109.870 -23.850 ;
        RECT 110.260 -24.280 110.670 -23.850 ;
        RECT 111.270 -23.920 111.720 -23.850 ;
        RECT 112.670 -23.610 113.120 -23.530 ;
        RECT 113.720 -23.610 114.130 -23.170 ;
        RECT 114.520 -23.610 114.970 -23.500 ;
        RECT 112.670 -23.850 114.970 -23.610 ;
        RECT 112.670 -23.950 113.120 -23.850 ;
        RECT 114.520 -23.950 114.970 -23.850 ;
        RECT 116.160 -23.610 116.610 -23.500 ;
        RECT 117.000 -23.610 117.410 -23.170 ;
        RECT 120.180 -23.440 120.630 -23.160 ;
        RECT 124.000 -23.440 124.450 -23.160 ;
        RECT 133.680 -23.160 135.210 -22.950 ;
        RECT 135.590 -23.040 136.040 -22.950 ;
        RECT 136.420 -23.160 137.950 -22.950 ;
        RECT 118.010 -23.610 118.460 -23.530 ;
        RECT 116.160 -23.850 118.460 -23.610 ;
        RECT 116.160 -23.950 116.610 -23.850 ;
        RECT 118.010 -23.950 118.460 -23.850 ;
        RECT 119.410 -23.610 119.860 -23.500 ;
        RECT 121.260 -23.610 121.710 -23.500 ;
        RECT 119.410 -23.850 121.710 -23.610 ;
        RECT 119.410 -23.920 119.860 -23.850 ;
        RECT 102.660 -24.480 103.110 -24.430 ;
        RECT 101.020 -24.770 103.110 -24.480 ;
        RECT 101.020 -24.820 101.470 -24.770 ;
        RECT 84.270 -25.400 84.720 -25.330 ;
        RECT 82.420 -25.640 84.720 -25.400 ;
        RECT 82.420 -25.750 82.870 -25.640 ;
        RECT 84.270 -25.750 84.720 -25.640 ;
        RECT 85.670 -25.400 86.120 -25.300 ;
        RECT 87.520 -25.400 87.970 -25.300 ;
        RECT 85.670 -25.640 87.970 -25.400 ;
        RECT 85.670 -25.720 86.120 -25.640 ;
        RECT 66.180 -26.300 67.710 -26.090 ;
        RECT 68.090 -26.300 68.540 -26.210 ;
        RECT 68.920 -26.300 70.450 -26.090 ;
        RECT 79.680 -26.090 80.130 -25.810 ;
        RECT 83.500 -26.090 83.950 -25.810 ;
        RECT 86.720 -26.080 87.130 -25.640 ;
        RECT 87.520 -25.750 87.970 -25.640 ;
        RECT 89.160 -25.400 89.610 -25.300 ;
        RECT 91.010 -25.400 91.460 -25.300 ;
        RECT 89.160 -25.640 91.460 -25.400 ;
        RECT 89.160 -25.750 89.610 -25.640 ;
        RECT 90.000 -26.080 90.410 -25.640 ;
        RECT 91.010 -25.720 91.460 -25.640 ;
        RECT 92.410 -25.400 92.860 -25.330 ;
        RECT 93.460 -25.400 93.870 -24.970 ;
        RECT 94.260 -25.400 94.710 -25.300 ;
        RECT 92.410 -25.640 94.710 -25.400 ;
        RECT 92.410 -25.750 92.860 -25.640 ;
        RECT 94.260 -25.750 94.710 -25.640 ;
        RECT 95.920 -25.400 96.370 -25.300 ;
        RECT 96.760 -25.400 97.170 -24.970 ;
        RECT 99.920 -25.040 101.470 -24.820 ;
        RECT 101.850 -24.830 102.280 -24.770 ;
        RECT 102.660 -24.820 103.110 -24.770 ;
        RECT 103.710 -24.820 104.210 -24.430 ;
        RECT 102.660 -25.040 104.210 -24.820 ;
        RECT 113.420 -24.430 114.970 -24.210 ;
        RECT 113.420 -24.820 113.920 -24.430 ;
        RECT 114.520 -24.480 114.970 -24.430 ;
        RECT 115.350 -24.480 115.780 -24.420 ;
        RECT 116.160 -24.430 117.710 -24.210 ;
        RECT 120.460 -24.280 120.870 -23.850 ;
        RECT 121.260 -23.950 121.710 -23.850 ;
        RECT 122.920 -23.610 123.370 -23.500 ;
        RECT 124.770 -23.610 125.220 -23.500 ;
        RECT 122.920 -23.850 125.220 -23.610 ;
        RECT 122.920 -23.950 123.370 -23.850 ;
        RECT 123.760 -24.280 124.170 -23.850 ;
        RECT 124.770 -23.920 125.220 -23.850 ;
        RECT 126.170 -23.610 126.620 -23.530 ;
        RECT 127.220 -23.610 127.630 -23.170 ;
        RECT 128.020 -23.610 128.470 -23.500 ;
        RECT 126.170 -23.850 128.470 -23.610 ;
        RECT 126.170 -23.950 126.620 -23.850 ;
        RECT 128.020 -23.950 128.470 -23.850 ;
        RECT 129.660 -23.610 130.110 -23.500 ;
        RECT 130.500 -23.610 130.910 -23.170 ;
        RECT 133.680 -23.440 134.130 -23.160 ;
        RECT 137.500 -23.440 137.950 -23.160 ;
        RECT 147.180 -23.160 148.710 -22.950 ;
        RECT 149.090 -23.040 149.540 -22.950 ;
        RECT 149.920 -23.160 151.450 -22.950 ;
        RECT 131.510 -23.610 131.960 -23.530 ;
        RECT 129.660 -23.850 131.960 -23.610 ;
        RECT 129.660 -23.950 130.110 -23.850 ;
        RECT 131.510 -23.950 131.960 -23.850 ;
        RECT 132.910 -23.610 133.360 -23.500 ;
        RECT 134.760 -23.610 135.210 -23.500 ;
        RECT 132.910 -23.850 135.210 -23.610 ;
        RECT 132.910 -23.920 133.360 -23.850 ;
        RECT 116.160 -24.480 116.610 -24.430 ;
        RECT 114.520 -24.770 116.610 -24.480 ;
        RECT 114.520 -24.820 114.970 -24.770 ;
        RECT 97.770 -25.400 98.220 -25.330 ;
        RECT 95.920 -25.640 98.220 -25.400 ;
        RECT 95.920 -25.750 96.370 -25.640 ;
        RECT 97.770 -25.750 98.220 -25.640 ;
        RECT 99.170 -25.400 99.620 -25.300 ;
        RECT 101.020 -25.400 101.470 -25.300 ;
        RECT 99.170 -25.640 101.470 -25.400 ;
        RECT 99.170 -25.720 99.620 -25.640 ;
        RECT 79.680 -26.300 81.210 -26.090 ;
        RECT 81.590 -26.300 82.040 -26.210 ;
        RECT 82.420 -26.300 83.950 -26.090 ;
        RECT 93.180 -26.090 93.630 -25.810 ;
        RECT 97.000 -26.090 97.450 -25.810 ;
        RECT 100.220 -26.080 100.630 -25.640 ;
        RECT 101.020 -25.750 101.470 -25.640 ;
        RECT 102.660 -25.400 103.110 -25.300 ;
        RECT 104.510 -25.400 104.960 -25.300 ;
        RECT 102.660 -25.640 104.960 -25.400 ;
        RECT 102.660 -25.750 103.110 -25.640 ;
        RECT 103.500 -26.080 103.910 -25.640 ;
        RECT 104.510 -25.720 104.960 -25.640 ;
        RECT 105.910 -25.400 106.360 -25.330 ;
        RECT 106.960 -25.400 107.370 -24.970 ;
        RECT 107.760 -25.400 108.210 -25.300 ;
        RECT 105.910 -25.640 108.210 -25.400 ;
        RECT 105.910 -25.750 106.360 -25.640 ;
        RECT 107.760 -25.750 108.210 -25.640 ;
        RECT 109.420 -25.400 109.870 -25.300 ;
        RECT 110.260 -25.400 110.670 -24.970 ;
        RECT 113.420 -25.040 114.970 -24.820 ;
        RECT 115.350 -24.830 115.780 -24.770 ;
        RECT 116.160 -24.820 116.610 -24.770 ;
        RECT 117.210 -24.820 117.710 -24.430 ;
        RECT 116.160 -25.040 117.710 -24.820 ;
        RECT 126.920 -24.430 128.470 -24.210 ;
        RECT 126.920 -24.820 127.420 -24.430 ;
        RECT 128.020 -24.480 128.470 -24.430 ;
        RECT 128.850 -24.480 129.280 -24.420 ;
        RECT 129.660 -24.430 131.210 -24.210 ;
        RECT 133.960 -24.280 134.370 -23.850 ;
        RECT 134.760 -23.950 135.210 -23.850 ;
        RECT 136.420 -23.610 136.870 -23.500 ;
        RECT 138.270 -23.610 138.720 -23.500 ;
        RECT 136.420 -23.850 138.720 -23.610 ;
        RECT 136.420 -23.950 136.870 -23.850 ;
        RECT 137.260 -24.280 137.670 -23.850 ;
        RECT 138.270 -23.920 138.720 -23.850 ;
        RECT 139.670 -23.610 140.120 -23.530 ;
        RECT 140.720 -23.610 141.130 -23.170 ;
        RECT 141.520 -23.610 141.970 -23.500 ;
        RECT 139.670 -23.850 141.970 -23.610 ;
        RECT 139.670 -23.950 140.120 -23.850 ;
        RECT 141.520 -23.950 141.970 -23.850 ;
        RECT 143.160 -23.610 143.610 -23.500 ;
        RECT 144.000 -23.610 144.410 -23.170 ;
        RECT 147.180 -23.440 147.630 -23.160 ;
        RECT 151.000 -23.440 151.450 -23.160 ;
        RECT 160.680 -23.160 162.210 -22.950 ;
        RECT 162.590 -23.040 163.040 -22.950 ;
        RECT 163.420 -23.160 164.950 -22.950 ;
        RECT 145.010 -23.610 145.460 -23.530 ;
        RECT 143.160 -23.850 145.460 -23.610 ;
        RECT 143.160 -23.950 143.610 -23.850 ;
        RECT 145.010 -23.950 145.460 -23.850 ;
        RECT 146.410 -23.610 146.860 -23.500 ;
        RECT 148.260 -23.610 148.710 -23.500 ;
        RECT 146.410 -23.850 148.710 -23.610 ;
        RECT 146.410 -23.920 146.860 -23.850 ;
        RECT 129.660 -24.480 130.110 -24.430 ;
        RECT 128.020 -24.770 130.110 -24.480 ;
        RECT 128.020 -24.820 128.470 -24.770 ;
        RECT 111.270 -25.400 111.720 -25.330 ;
        RECT 109.420 -25.640 111.720 -25.400 ;
        RECT 109.420 -25.750 109.870 -25.640 ;
        RECT 111.270 -25.750 111.720 -25.640 ;
        RECT 112.670 -25.400 113.120 -25.300 ;
        RECT 114.520 -25.400 114.970 -25.300 ;
        RECT 112.670 -25.640 114.970 -25.400 ;
        RECT 112.670 -25.720 113.120 -25.640 ;
        RECT 93.180 -26.300 94.710 -26.090 ;
        RECT 95.090 -26.300 95.540 -26.210 ;
        RECT 95.920 -26.300 97.450 -26.090 ;
        RECT 106.680 -26.090 107.130 -25.810 ;
        RECT 110.500 -26.090 110.950 -25.810 ;
        RECT 113.720 -26.080 114.130 -25.640 ;
        RECT 114.520 -25.750 114.970 -25.640 ;
        RECT 116.160 -25.400 116.610 -25.300 ;
        RECT 118.010 -25.400 118.460 -25.300 ;
        RECT 116.160 -25.640 118.460 -25.400 ;
        RECT 116.160 -25.750 116.610 -25.640 ;
        RECT 117.000 -26.080 117.410 -25.640 ;
        RECT 118.010 -25.720 118.460 -25.640 ;
        RECT 119.410 -25.400 119.860 -25.330 ;
        RECT 120.460 -25.400 120.870 -24.970 ;
        RECT 121.260 -25.400 121.710 -25.300 ;
        RECT 119.410 -25.640 121.710 -25.400 ;
        RECT 119.410 -25.750 119.860 -25.640 ;
        RECT 121.260 -25.750 121.710 -25.640 ;
        RECT 122.920 -25.400 123.370 -25.300 ;
        RECT 123.760 -25.400 124.170 -24.970 ;
        RECT 126.920 -25.040 128.470 -24.820 ;
        RECT 128.850 -24.830 129.280 -24.770 ;
        RECT 129.660 -24.820 130.110 -24.770 ;
        RECT 130.710 -24.820 131.210 -24.430 ;
        RECT 129.660 -25.040 131.210 -24.820 ;
        RECT 140.420 -24.430 141.970 -24.210 ;
        RECT 140.420 -24.820 140.920 -24.430 ;
        RECT 141.520 -24.480 141.970 -24.430 ;
        RECT 142.350 -24.480 142.780 -24.420 ;
        RECT 143.160 -24.430 144.710 -24.210 ;
        RECT 147.460 -24.280 147.870 -23.850 ;
        RECT 148.260 -23.950 148.710 -23.850 ;
        RECT 149.920 -23.610 150.370 -23.500 ;
        RECT 151.770 -23.610 152.220 -23.500 ;
        RECT 149.920 -23.850 152.220 -23.610 ;
        RECT 149.920 -23.950 150.370 -23.850 ;
        RECT 150.760 -24.280 151.170 -23.850 ;
        RECT 151.770 -23.920 152.220 -23.850 ;
        RECT 153.170 -23.610 153.620 -23.530 ;
        RECT 154.220 -23.610 154.630 -23.170 ;
        RECT 155.020 -23.610 155.470 -23.500 ;
        RECT 153.170 -23.850 155.470 -23.610 ;
        RECT 153.170 -23.950 153.620 -23.850 ;
        RECT 155.020 -23.950 155.470 -23.850 ;
        RECT 156.660 -23.610 157.110 -23.500 ;
        RECT 157.500 -23.610 157.910 -23.170 ;
        RECT 160.680 -23.440 161.130 -23.160 ;
        RECT 164.500 -23.440 164.950 -23.160 ;
        RECT 174.180 -23.160 175.710 -22.950 ;
        RECT 176.090 -23.040 176.540 -22.950 ;
        RECT 176.920 -23.160 178.450 -22.950 ;
        RECT 158.510 -23.610 158.960 -23.530 ;
        RECT 156.660 -23.850 158.960 -23.610 ;
        RECT 156.660 -23.950 157.110 -23.850 ;
        RECT 158.510 -23.950 158.960 -23.850 ;
        RECT 159.910 -23.610 160.360 -23.500 ;
        RECT 161.760 -23.610 162.210 -23.500 ;
        RECT 159.910 -23.850 162.210 -23.610 ;
        RECT 159.910 -23.920 160.360 -23.850 ;
        RECT 143.160 -24.480 143.610 -24.430 ;
        RECT 141.520 -24.770 143.610 -24.480 ;
        RECT 141.520 -24.820 141.970 -24.770 ;
        RECT 124.770 -25.400 125.220 -25.330 ;
        RECT 122.920 -25.640 125.220 -25.400 ;
        RECT 122.920 -25.750 123.370 -25.640 ;
        RECT 124.770 -25.750 125.220 -25.640 ;
        RECT 126.170 -25.400 126.620 -25.300 ;
        RECT 128.020 -25.400 128.470 -25.300 ;
        RECT 126.170 -25.640 128.470 -25.400 ;
        RECT 126.170 -25.720 126.620 -25.640 ;
        RECT 106.680 -26.250 108.210 -26.090 ;
        RECT 108.590 -26.250 109.040 -26.210 ;
        RECT 109.420 -26.250 110.950 -26.090 ;
        RECT 106.680 -26.300 110.950 -26.250 ;
        RECT 120.180 -26.090 120.630 -25.810 ;
        RECT 124.000 -26.090 124.450 -25.810 ;
        RECT 127.220 -26.080 127.630 -25.640 ;
        RECT 128.020 -25.750 128.470 -25.640 ;
        RECT 129.660 -25.400 130.110 -25.300 ;
        RECT 131.510 -25.400 131.960 -25.300 ;
        RECT 129.660 -25.640 131.960 -25.400 ;
        RECT 129.660 -25.750 130.110 -25.640 ;
        RECT 130.500 -26.080 130.910 -25.640 ;
        RECT 131.510 -25.720 131.960 -25.640 ;
        RECT 132.910 -25.400 133.360 -25.330 ;
        RECT 133.960 -25.400 134.370 -24.970 ;
        RECT 134.760 -25.400 135.210 -25.300 ;
        RECT 132.910 -25.640 135.210 -25.400 ;
        RECT 132.910 -25.750 133.360 -25.640 ;
        RECT 134.760 -25.750 135.210 -25.640 ;
        RECT 136.420 -25.400 136.870 -25.300 ;
        RECT 137.260 -25.400 137.670 -24.970 ;
        RECT 140.420 -25.040 141.970 -24.820 ;
        RECT 142.350 -24.830 142.780 -24.770 ;
        RECT 143.160 -24.820 143.610 -24.770 ;
        RECT 144.210 -24.820 144.710 -24.430 ;
        RECT 143.160 -25.040 144.710 -24.820 ;
        RECT 153.920 -24.430 155.470 -24.210 ;
        RECT 153.920 -24.820 154.420 -24.430 ;
        RECT 155.020 -24.480 155.470 -24.430 ;
        RECT 155.850 -24.480 156.280 -24.420 ;
        RECT 156.660 -24.430 158.210 -24.210 ;
        RECT 160.960 -24.280 161.370 -23.850 ;
        RECT 161.760 -23.950 162.210 -23.850 ;
        RECT 163.420 -23.610 163.870 -23.500 ;
        RECT 165.270 -23.610 165.720 -23.500 ;
        RECT 163.420 -23.850 165.720 -23.610 ;
        RECT 163.420 -23.950 163.870 -23.850 ;
        RECT 164.260 -24.280 164.670 -23.850 ;
        RECT 165.270 -23.920 165.720 -23.850 ;
        RECT 166.670 -23.610 167.120 -23.530 ;
        RECT 167.720 -23.610 168.130 -23.170 ;
        RECT 168.520 -23.610 168.970 -23.500 ;
        RECT 166.670 -23.850 168.970 -23.610 ;
        RECT 166.670 -23.950 167.120 -23.850 ;
        RECT 168.520 -23.950 168.970 -23.850 ;
        RECT 170.160 -23.610 170.610 -23.500 ;
        RECT 171.000 -23.610 171.410 -23.170 ;
        RECT 174.180 -23.440 174.630 -23.160 ;
        RECT 178.000 -23.440 178.450 -23.160 ;
        RECT 187.680 -23.160 189.210 -22.950 ;
        RECT 189.590 -23.040 190.040 -22.950 ;
        RECT 190.420 -23.160 191.950 -22.950 ;
        RECT 172.010 -23.610 172.460 -23.530 ;
        RECT 170.160 -23.850 172.460 -23.610 ;
        RECT 170.160 -23.950 170.610 -23.850 ;
        RECT 172.010 -23.950 172.460 -23.850 ;
        RECT 173.410 -23.610 173.860 -23.500 ;
        RECT 175.260 -23.610 175.710 -23.500 ;
        RECT 173.410 -23.850 175.710 -23.610 ;
        RECT 173.410 -23.920 173.860 -23.850 ;
        RECT 156.660 -24.480 157.110 -24.430 ;
        RECT 155.020 -24.770 157.110 -24.480 ;
        RECT 155.020 -24.820 155.470 -24.770 ;
        RECT 138.270 -25.400 138.720 -25.330 ;
        RECT 136.420 -25.640 138.720 -25.400 ;
        RECT 136.420 -25.750 136.870 -25.640 ;
        RECT 138.270 -25.750 138.720 -25.640 ;
        RECT 139.670 -25.400 140.120 -25.300 ;
        RECT 141.520 -25.400 141.970 -25.300 ;
        RECT 139.670 -25.640 141.970 -25.400 ;
        RECT 139.670 -25.720 140.120 -25.640 ;
        RECT 120.180 -26.300 121.710 -26.090 ;
        RECT 122.090 -26.300 122.540 -26.210 ;
        RECT 122.920 -26.300 124.450 -26.090 ;
        RECT 133.680 -26.090 134.130 -25.810 ;
        RECT 137.500 -26.090 137.950 -25.810 ;
        RECT 140.720 -26.080 141.130 -25.640 ;
        RECT 141.520 -25.750 141.970 -25.640 ;
        RECT 143.160 -25.400 143.610 -25.300 ;
        RECT 145.010 -25.400 145.460 -25.300 ;
        RECT 143.160 -25.640 145.460 -25.400 ;
        RECT 143.160 -25.750 143.610 -25.640 ;
        RECT 144.000 -26.080 144.410 -25.640 ;
        RECT 145.010 -25.720 145.460 -25.640 ;
        RECT 146.410 -25.400 146.860 -25.330 ;
        RECT 147.460 -25.400 147.870 -24.970 ;
        RECT 148.260 -25.400 148.710 -25.300 ;
        RECT 146.410 -25.640 148.710 -25.400 ;
        RECT 146.410 -25.750 146.860 -25.640 ;
        RECT 148.260 -25.750 148.710 -25.640 ;
        RECT 149.920 -25.400 150.370 -25.300 ;
        RECT 150.760 -25.400 151.170 -24.970 ;
        RECT 153.920 -25.040 155.470 -24.820 ;
        RECT 155.850 -24.830 156.280 -24.770 ;
        RECT 156.660 -24.820 157.110 -24.770 ;
        RECT 157.710 -24.820 158.210 -24.430 ;
        RECT 156.660 -25.040 158.210 -24.820 ;
        RECT 167.420 -24.430 168.970 -24.210 ;
        RECT 167.420 -24.820 167.920 -24.430 ;
        RECT 168.520 -24.480 168.970 -24.430 ;
        RECT 169.350 -24.480 169.780 -24.420 ;
        RECT 170.160 -24.430 171.710 -24.210 ;
        RECT 174.460 -24.280 174.870 -23.850 ;
        RECT 175.260 -23.950 175.710 -23.850 ;
        RECT 176.920 -23.610 177.370 -23.500 ;
        RECT 178.770 -23.610 179.220 -23.500 ;
        RECT 176.920 -23.850 179.220 -23.610 ;
        RECT 176.920 -23.950 177.370 -23.850 ;
        RECT 177.760 -24.280 178.170 -23.850 ;
        RECT 178.770 -23.920 179.220 -23.850 ;
        RECT 180.170 -23.610 180.620 -23.530 ;
        RECT 181.220 -23.610 181.630 -23.170 ;
        RECT 182.020 -23.610 182.470 -23.500 ;
        RECT 180.170 -23.850 182.470 -23.610 ;
        RECT 180.170 -23.950 180.620 -23.850 ;
        RECT 182.020 -23.950 182.470 -23.850 ;
        RECT 183.660 -23.610 184.110 -23.500 ;
        RECT 184.500 -23.610 184.910 -23.170 ;
        RECT 187.680 -23.440 188.130 -23.160 ;
        RECT 191.500 -23.440 191.950 -23.160 ;
        RECT 201.180 -23.160 202.710 -22.950 ;
        RECT 203.090 -23.040 203.540 -22.950 ;
        RECT 203.920 -23.160 205.450 -22.950 ;
        RECT 185.510 -23.610 185.960 -23.530 ;
        RECT 183.660 -23.850 185.960 -23.610 ;
        RECT 183.660 -23.950 184.110 -23.850 ;
        RECT 185.510 -23.950 185.960 -23.850 ;
        RECT 186.910 -23.610 187.360 -23.500 ;
        RECT 188.760 -23.610 189.210 -23.500 ;
        RECT 186.910 -23.850 189.210 -23.610 ;
        RECT 186.910 -23.920 187.360 -23.850 ;
        RECT 170.160 -24.480 170.610 -24.430 ;
        RECT 168.520 -24.770 170.610 -24.480 ;
        RECT 168.520 -24.820 168.970 -24.770 ;
        RECT 151.770 -25.400 152.220 -25.330 ;
        RECT 149.920 -25.640 152.220 -25.400 ;
        RECT 149.920 -25.750 150.370 -25.640 ;
        RECT 151.770 -25.750 152.220 -25.640 ;
        RECT 153.170 -25.400 153.620 -25.300 ;
        RECT 155.020 -25.400 155.470 -25.300 ;
        RECT 153.170 -25.640 155.470 -25.400 ;
        RECT 153.170 -25.720 153.620 -25.640 ;
        RECT 133.680 -26.300 135.210 -26.090 ;
        RECT 135.590 -26.300 136.040 -26.210 ;
        RECT 136.420 -26.300 137.950 -26.090 ;
        RECT 147.180 -26.090 147.630 -25.810 ;
        RECT 151.000 -26.090 151.450 -25.810 ;
        RECT 154.220 -26.080 154.630 -25.640 ;
        RECT 155.020 -25.750 155.470 -25.640 ;
        RECT 156.660 -25.400 157.110 -25.300 ;
        RECT 158.510 -25.400 158.960 -25.300 ;
        RECT 156.660 -25.640 158.960 -25.400 ;
        RECT 156.660 -25.750 157.110 -25.640 ;
        RECT 157.500 -26.080 157.910 -25.640 ;
        RECT 158.510 -25.720 158.960 -25.640 ;
        RECT 159.910 -25.400 160.360 -25.330 ;
        RECT 160.960 -25.400 161.370 -24.970 ;
        RECT 161.760 -25.400 162.210 -25.300 ;
        RECT 159.910 -25.640 162.210 -25.400 ;
        RECT 159.910 -25.750 160.360 -25.640 ;
        RECT 161.760 -25.750 162.210 -25.640 ;
        RECT 163.420 -25.400 163.870 -25.300 ;
        RECT 164.260 -25.400 164.670 -24.970 ;
        RECT 167.420 -25.040 168.970 -24.820 ;
        RECT 169.350 -24.830 169.780 -24.770 ;
        RECT 170.160 -24.820 170.610 -24.770 ;
        RECT 171.210 -24.820 171.710 -24.430 ;
        RECT 170.160 -25.040 171.710 -24.820 ;
        RECT 180.920 -24.430 182.470 -24.210 ;
        RECT 180.920 -24.820 181.420 -24.430 ;
        RECT 182.020 -24.480 182.470 -24.430 ;
        RECT 182.850 -24.480 183.280 -24.420 ;
        RECT 183.660 -24.430 185.210 -24.210 ;
        RECT 187.960 -24.280 188.370 -23.850 ;
        RECT 188.760 -23.950 189.210 -23.850 ;
        RECT 190.420 -23.610 190.870 -23.500 ;
        RECT 192.270 -23.610 192.720 -23.500 ;
        RECT 190.420 -23.850 192.720 -23.610 ;
        RECT 190.420 -23.950 190.870 -23.850 ;
        RECT 191.260 -24.280 191.670 -23.850 ;
        RECT 192.270 -23.920 192.720 -23.850 ;
        RECT 193.670 -23.610 194.120 -23.530 ;
        RECT 194.720 -23.610 195.130 -23.170 ;
        RECT 195.520 -23.610 195.970 -23.500 ;
        RECT 193.670 -23.850 195.970 -23.610 ;
        RECT 193.670 -23.950 194.120 -23.850 ;
        RECT 195.520 -23.950 195.970 -23.850 ;
        RECT 197.160 -23.610 197.610 -23.500 ;
        RECT 198.000 -23.610 198.410 -23.170 ;
        RECT 201.180 -23.440 201.630 -23.160 ;
        RECT 205.000 -23.440 205.450 -23.160 ;
        RECT 214.680 -23.160 216.210 -22.950 ;
        RECT 216.590 -23.040 217.030 -22.950 ;
        RECT 199.010 -23.610 199.460 -23.530 ;
        RECT 197.160 -23.850 199.460 -23.610 ;
        RECT 197.160 -23.950 197.610 -23.850 ;
        RECT 199.010 -23.950 199.460 -23.850 ;
        RECT 200.410 -23.610 200.860 -23.500 ;
        RECT 202.260 -23.610 202.710 -23.500 ;
        RECT 200.410 -23.850 202.710 -23.610 ;
        RECT 200.410 -23.920 200.860 -23.850 ;
        RECT 183.660 -24.480 184.110 -24.430 ;
        RECT 182.020 -24.770 184.110 -24.480 ;
        RECT 182.020 -24.820 182.470 -24.770 ;
        RECT 165.270 -25.400 165.720 -25.330 ;
        RECT 163.420 -25.640 165.720 -25.400 ;
        RECT 163.420 -25.750 163.870 -25.640 ;
        RECT 165.270 -25.750 165.720 -25.640 ;
        RECT 166.670 -25.400 167.120 -25.300 ;
        RECT 168.520 -25.400 168.970 -25.300 ;
        RECT 166.670 -25.640 168.970 -25.400 ;
        RECT 166.670 -25.720 167.120 -25.640 ;
        RECT 147.180 -26.300 148.710 -26.090 ;
        RECT 149.090 -26.300 149.540 -26.210 ;
        RECT 149.920 -26.300 151.450 -26.090 ;
        RECT 160.680 -26.090 161.130 -25.810 ;
        RECT 164.500 -26.090 164.950 -25.810 ;
        RECT 167.720 -26.080 168.130 -25.640 ;
        RECT 168.520 -25.750 168.970 -25.640 ;
        RECT 170.160 -25.400 170.610 -25.300 ;
        RECT 172.010 -25.400 172.460 -25.300 ;
        RECT 170.160 -25.640 172.460 -25.400 ;
        RECT 170.160 -25.750 170.610 -25.640 ;
        RECT 171.000 -26.080 171.410 -25.640 ;
        RECT 172.010 -25.720 172.460 -25.640 ;
        RECT 173.410 -25.400 173.860 -25.330 ;
        RECT 174.460 -25.400 174.870 -24.970 ;
        RECT 175.260 -25.400 175.710 -25.300 ;
        RECT 173.410 -25.640 175.710 -25.400 ;
        RECT 173.410 -25.750 173.860 -25.640 ;
        RECT 175.260 -25.750 175.710 -25.640 ;
        RECT 176.920 -25.400 177.370 -25.300 ;
        RECT 177.760 -25.400 178.170 -24.970 ;
        RECT 180.920 -25.040 182.470 -24.820 ;
        RECT 182.850 -24.830 183.280 -24.770 ;
        RECT 183.660 -24.820 184.110 -24.770 ;
        RECT 184.710 -24.820 185.210 -24.430 ;
        RECT 183.660 -25.040 185.210 -24.820 ;
        RECT 194.420 -24.430 195.970 -24.210 ;
        RECT 194.420 -24.820 194.920 -24.430 ;
        RECT 195.520 -24.480 195.970 -24.430 ;
        RECT 196.350 -24.480 196.780 -24.420 ;
        RECT 197.160 -24.430 198.710 -24.210 ;
        RECT 201.460 -24.280 201.870 -23.850 ;
        RECT 202.260 -23.950 202.710 -23.850 ;
        RECT 203.920 -23.610 204.370 -23.500 ;
        RECT 205.770 -23.610 206.220 -23.500 ;
        RECT 203.920 -23.850 206.220 -23.610 ;
        RECT 203.920 -23.950 204.370 -23.850 ;
        RECT 204.760 -24.280 205.170 -23.850 ;
        RECT 205.770 -23.920 206.220 -23.850 ;
        RECT 207.170 -23.610 207.620 -23.530 ;
        RECT 208.220 -23.610 208.630 -23.170 ;
        RECT 209.020 -23.610 209.470 -23.500 ;
        RECT 207.170 -23.850 209.470 -23.610 ;
        RECT 207.170 -23.950 207.620 -23.850 ;
        RECT 209.020 -23.950 209.470 -23.850 ;
        RECT 210.660 -23.610 211.110 -23.500 ;
        RECT 211.500 -23.610 211.910 -23.170 ;
        RECT 214.680 -23.440 215.130 -23.160 ;
        RECT 212.510 -23.610 212.960 -23.530 ;
        RECT 210.660 -23.850 212.960 -23.610 ;
        RECT 210.660 -23.950 211.110 -23.850 ;
        RECT 212.510 -23.950 212.960 -23.850 ;
        RECT 213.910 -23.610 214.360 -23.500 ;
        RECT 215.760 -23.610 216.210 -23.500 ;
        RECT 213.910 -23.850 216.210 -23.610 ;
        RECT 213.910 -23.920 214.360 -23.850 ;
        RECT 197.160 -24.480 197.610 -24.430 ;
        RECT 195.520 -24.770 197.610 -24.480 ;
        RECT 195.520 -24.820 195.970 -24.770 ;
        RECT 178.770 -25.400 179.220 -25.330 ;
        RECT 176.920 -25.640 179.220 -25.400 ;
        RECT 176.920 -25.750 177.370 -25.640 ;
        RECT 178.770 -25.750 179.220 -25.640 ;
        RECT 180.170 -25.400 180.620 -25.300 ;
        RECT 182.020 -25.400 182.470 -25.300 ;
        RECT 180.170 -25.640 182.470 -25.400 ;
        RECT 180.170 -25.720 180.620 -25.640 ;
        RECT 160.680 -26.250 162.210 -26.090 ;
        RECT 162.590 -26.250 163.040 -26.210 ;
        RECT 163.420 -26.250 164.950 -26.090 ;
        RECT 160.680 -26.300 164.950 -26.250 ;
        RECT 174.180 -26.090 174.630 -25.810 ;
        RECT 178.000 -26.090 178.450 -25.810 ;
        RECT 181.220 -26.080 181.630 -25.640 ;
        RECT 182.020 -25.750 182.470 -25.640 ;
        RECT 183.660 -25.400 184.110 -25.300 ;
        RECT 185.510 -25.400 185.960 -25.300 ;
        RECT 183.660 -25.640 185.960 -25.400 ;
        RECT 183.660 -25.750 184.110 -25.640 ;
        RECT 184.500 -26.080 184.910 -25.640 ;
        RECT 185.510 -25.720 185.960 -25.640 ;
        RECT 186.910 -25.400 187.360 -25.330 ;
        RECT 187.960 -25.400 188.370 -24.970 ;
        RECT 188.760 -25.400 189.210 -25.300 ;
        RECT 186.910 -25.640 189.210 -25.400 ;
        RECT 186.910 -25.750 187.360 -25.640 ;
        RECT 188.760 -25.750 189.210 -25.640 ;
        RECT 190.420 -25.400 190.870 -25.300 ;
        RECT 191.260 -25.400 191.670 -24.970 ;
        RECT 194.420 -25.040 195.970 -24.820 ;
        RECT 196.350 -24.830 196.780 -24.770 ;
        RECT 197.160 -24.820 197.610 -24.770 ;
        RECT 198.210 -24.820 198.710 -24.430 ;
        RECT 197.160 -25.040 198.710 -24.820 ;
        RECT 207.920 -24.430 209.470 -24.210 ;
        RECT 207.920 -24.820 208.420 -24.430 ;
        RECT 209.020 -24.480 209.470 -24.430 ;
        RECT 209.850 -24.480 210.280 -24.420 ;
        RECT 210.660 -24.430 212.210 -24.210 ;
        RECT 214.960 -24.280 215.370 -23.850 ;
        RECT 215.760 -23.950 216.210 -23.850 ;
        RECT 210.660 -24.480 211.110 -24.430 ;
        RECT 209.020 -24.770 211.110 -24.480 ;
        RECT 209.020 -24.820 209.470 -24.770 ;
        RECT 192.270 -25.400 192.720 -25.330 ;
        RECT 190.420 -25.640 192.720 -25.400 ;
        RECT 190.420 -25.750 190.870 -25.640 ;
        RECT 192.270 -25.750 192.720 -25.640 ;
        RECT 193.670 -25.400 194.120 -25.300 ;
        RECT 195.520 -25.400 195.970 -25.300 ;
        RECT 193.670 -25.640 195.970 -25.400 ;
        RECT 193.670 -25.720 194.120 -25.640 ;
        RECT 174.180 -26.300 175.710 -26.090 ;
        RECT 176.090 -26.300 176.540 -26.210 ;
        RECT 176.920 -26.300 178.450 -26.090 ;
        RECT 187.680 -26.090 188.130 -25.810 ;
        RECT 191.500 -26.090 191.950 -25.810 ;
        RECT 194.720 -26.080 195.130 -25.640 ;
        RECT 195.520 -25.750 195.970 -25.640 ;
        RECT 197.160 -25.400 197.610 -25.300 ;
        RECT 199.010 -25.400 199.460 -25.300 ;
        RECT 197.160 -25.640 199.460 -25.400 ;
        RECT 197.160 -25.750 197.610 -25.640 ;
        RECT 198.000 -26.080 198.410 -25.640 ;
        RECT 199.010 -25.720 199.460 -25.640 ;
        RECT 200.410 -25.400 200.860 -25.330 ;
        RECT 201.460 -25.400 201.870 -24.970 ;
        RECT 202.260 -25.400 202.710 -25.300 ;
        RECT 200.410 -25.640 202.710 -25.400 ;
        RECT 200.410 -25.750 200.860 -25.640 ;
        RECT 202.260 -25.750 202.710 -25.640 ;
        RECT 203.920 -25.400 204.370 -25.300 ;
        RECT 204.760 -25.400 205.170 -24.970 ;
        RECT 207.920 -25.040 209.470 -24.820 ;
        RECT 209.850 -24.830 210.280 -24.770 ;
        RECT 210.660 -24.820 211.110 -24.770 ;
        RECT 211.710 -24.820 212.210 -24.430 ;
        RECT 210.660 -25.040 212.210 -24.820 ;
        RECT 205.770 -25.400 206.220 -25.330 ;
        RECT 203.920 -25.640 206.220 -25.400 ;
        RECT 203.920 -25.750 204.370 -25.640 ;
        RECT 205.770 -25.750 206.220 -25.640 ;
        RECT 207.170 -25.400 207.620 -25.300 ;
        RECT 209.020 -25.400 209.470 -25.300 ;
        RECT 207.170 -25.640 209.470 -25.400 ;
        RECT 207.170 -25.720 207.620 -25.640 ;
        RECT 187.680 -26.300 189.210 -26.090 ;
        RECT 189.590 -26.300 190.040 -26.210 ;
        RECT 190.420 -26.300 191.950 -26.090 ;
        RECT 201.180 -26.090 201.630 -25.810 ;
        RECT 205.000 -26.090 205.450 -25.810 ;
        RECT 208.220 -26.080 208.630 -25.640 ;
        RECT 209.020 -25.750 209.470 -25.640 ;
        RECT 210.660 -25.400 211.110 -25.300 ;
        RECT 212.510 -25.400 212.960 -25.300 ;
        RECT 210.660 -25.640 212.960 -25.400 ;
        RECT 210.660 -25.750 211.110 -25.640 ;
        RECT 211.500 -26.080 211.910 -25.640 ;
        RECT 212.510 -25.720 212.960 -25.640 ;
        RECT 213.910 -25.400 214.360 -25.330 ;
        RECT 214.960 -25.400 215.370 -24.970 ;
        RECT 215.760 -25.400 216.210 -25.300 ;
        RECT 213.910 -25.640 216.210 -25.400 ;
        RECT 213.910 -25.750 214.360 -25.640 ;
        RECT 215.760 -25.750 216.210 -25.640 ;
        RECT 201.180 -26.300 202.710 -26.090 ;
        RECT 203.090 -26.300 203.540 -26.210 ;
        RECT 203.920 -26.300 205.450 -26.090 ;
        RECT 214.680 -26.090 215.130 -25.810 ;
        RECT 214.680 -26.300 216.210 -26.090 ;
        RECT 216.590 -26.250 217.030 -26.210 ;
        RECT 216.590 -26.300 217.690 -26.250 ;
        RECT 13.260 -26.560 15.370 -26.300 ;
        RECT 26.760 -26.560 28.870 -26.300 ;
        RECT 40.260 -26.560 42.370 -26.300 ;
        RECT 53.760 -26.560 55.870 -26.300 ;
        RECT 67.260 -26.560 69.370 -26.300 ;
        RECT 80.760 -26.560 82.870 -26.300 ;
        RECT 94.260 -26.560 96.370 -26.300 ;
        RECT 107.760 -26.560 109.870 -26.300 ;
        RECT 121.260 -26.560 123.370 -26.300 ;
        RECT 134.760 -26.560 136.870 -26.300 ;
        RECT 148.260 -26.560 150.370 -26.300 ;
        RECT 161.760 -26.560 163.870 -26.300 ;
        RECT 175.260 -26.560 177.370 -26.300 ;
        RECT 188.760 -26.560 190.870 -26.300 ;
        RECT 202.260 -26.560 204.370 -26.300 ;
        RECT 215.760 -26.560 217.690 -26.300 ;
        RECT 12.180 -26.770 13.710 -26.560 ;
        RECT 14.090 -26.650 14.540 -26.560 ;
        RECT 14.920 -26.770 16.450 -26.560 ;
        RECT 1.420 -27.220 1.870 -27.110 ;
        RECT 3.270 -27.220 3.720 -27.110 ;
        RECT 1.420 -27.460 3.720 -27.220 ;
        RECT 1.420 -27.560 1.870 -27.460 ;
        RECT 2.260 -27.890 2.670 -27.460 ;
        RECT 3.270 -27.530 3.720 -27.460 ;
        RECT 4.670 -27.220 5.120 -27.140 ;
        RECT 5.720 -27.220 6.130 -26.780 ;
        RECT 6.520 -27.220 6.970 -27.110 ;
        RECT 4.670 -27.460 6.970 -27.220 ;
        RECT 4.670 -27.560 5.120 -27.460 ;
        RECT 6.520 -27.560 6.970 -27.460 ;
        RECT 8.160 -27.220 8.610 -27.110 ;
        RECT 9.000 -27.220 9.410 -26.780 ;
        RECT 12.180 -27.050 12.630 -26.770 ;
        RECT 16.000 -27.050 16.450 -26.770 ;
        RECT 25.680 -26.770 27.210 -26.560 ;
        RECT 27.590 -26.650 28.040 -26.560 ;
        RECT 28.420 -26.770 29.950 -26.560 ;
        RECT 10.010 -27.220 10.460 -27.140 ;
        RECT 8.160 -27.460 10.460 -27.220 ;
        RECT 8.160 -27.560 8.610 -27.460 ;
        RECT 10.010 -27.560 10.460 -27.460 ;
        RECT 11.410 -27.220 11.860 -27.110 ;
        RECT 13.260 -27.220 13.710 -27.110 ;
        RECT 11.410 -27.460 13.710 -27.220 ;
        RECT 11.410 -27.530 11.860 -27.460 ;
        RECT 5.420 -28.040 6.970 -27.820 ;
        RECT 5.420 -28.430 5.920 -28.040 ;
        RECT 6.520 -28.090 6.970 -28.040 ;
        RECT 7.350 -28.090 7.780 -28.030 ;
        RECT 8.160 -28.040 9.710 -27.820 ;
        RECT 12.460 -27.890 12.870 -27.460 ;
        RECT 13.260 -27.560 13.710 -27.460 ;
        RECT 14.920 -27.220 15.370 -27.110 ;
        RECT 16.770 -27.220 17.220 -27.110 ;
        RECT 14.920 -27.460 17.220 -27.220 ;
        RECT 14.920 -27.560 15.370 -27.460 ;
        RECT 15.760 -27.890 16.170 -27.460 ;
        RECT 16.770 -27.530 17.220 -27.460 ;
        RECT 18.170 -27.220 18.620 -27.140 ;
        RECT 19.220 -27.220 19.630 -26.780 ;
        RECT 20.020 -27.220 20.470 -27.110 ;
        RECT 18.170 -27.460 20.470 -27.220 ;
        RECT 18.170 -27.560 18.620 -27.460 ;
        RECT 20.020 -27.560 20.470 -27.460 ;
        RECT 21.660 -27.220 22.110 -27.110 ;
        RECT 22.500 -27.220 22.910 -26.780 ;
        RECT 25.680 -27.050 26.130 -26.770 ;
        RECT 29.500 -27.050 29.950 -26.770 ;
        RECT 39.180 -26.770 40.710 -26.560 ;
        RECT 41.090 -26.650 41.540 -26.560 ;
        RECT 41.920 -26.770 43.450 -26.560 ;
        RECT 23.510 -27.220 23.960 -27.140 ;
        RECT 21.660 -27.460 23.960 -27.220 ;
        RECT 21.660 -27.560 22.110 -27.460 ;
        RECT 23.510 -27.560 23.960 -27.460 ;
        RECT 24.910 -27.220 25.360 -27.110 ;
        RECT 26.760 -27.220 27.210 -27.110 ;
        RECT 24.910 -27.460 27.210 -27.220 ;
        RECT 24.910 -27.530 25.360 -27.460 ;
        RECT 8.160 -28.090 8.610 -28.040 ;
        RECT 6.520 -28.380 8.610 -28.090 ;
        RECT 6.520 -28.430 6.970 -28.380 ;
        RECT 1.420 -29.010 1.870 -28.910 ;
        RECT 2.260 -29.010 2.670 -28.580 ;
        RECT 5.420 -28.650 6.970 -28.430 ;
        RECT 7.350 -28.440 7.780 -28.380 ;
        RECT 8.160 -28.430 8.610 -28.380 ;
        RECT 9.210 -28.430 9.710 -28.040 ;
        RECT 8.160 -28.650 9.710 -28.430 ;
        RECT 18.920 -28.040 20.470 -27.820 ;
        RECT 18.920 -28.430 19.420 -28.040 ;
        RECT 20.020 -28.090 20.470 -28.040 ;
        RECT 20.850 -28.090 21.280 -28.030 ;
        RECT 21.660 -28.040 23.210 -27.820 ;
        RECT 25.960 -27.890 26.370 -27.460 ;
        RECT 26.760 -27.560 27.210 -27.460 ;
        RECT 28.420 -27.220 28.870 -27.110 ;
        RECT 30.270 -27.220 30.720 -27.110 ;
        RECT 28.420 -27.460 30.720 -27.220 ;
        RECT 28.420 -27.560 28.870 -27.460 ;
        RECT 29.260 -27.890 29.670 -27.460 ;
        RECT 30.270 -27.530 30.720 -27.460 ;
        RECT 31.670 -27.220 32.120 -27.140 ;
        RECT 32.720 -27.220 33.130 -26.780 ;
        RECT 33.520 -27.220 33.970 -27.110 ;
        RECT 31.670 -27.460 33.970 -27.220 ;
        RECT 31.670 -27.560 32.120 -27.460 ;
        RECT 33.520 -27.560 33.970 -27.460 ;
        RECT 35.160 -27.220 35.610 -27.110 ;
        RECT 36.000 -27.220 36.410 -26.780 ;
        RECT 39.180 -27.050 39.630 -26.770 ;
        RECT 43.000 -27.050 43.450 -26.770 ;
        RECT 52.680 -26.610 56.950 -26.560 ;
        RECT 52.680 -26.770 54.210 -26.610 ;
        RECT 54.590 -26.650 55.040 -26.610 ;
        RECT 55.420 -26.770 56.950 -26.610 ;
        RECT 37.010 -27.220 37.460 -27.140 ;
        RECT 35.160 -27.460 37.460 -27.220 ;
        RECT 35.160 -27.560 35.610 -27.460 ;
        RECT 37.010 -27.560 37.460 -27.460 ;
        RECT 38.410 -27.220 38.860 -27.110 ;
        RECT 40.260 -27.220 40.710 -27.110 ;
        RECT 38.410 -27.460 40.710 -27.220 ;
        RECT 38.410 -27.530 38.860 -27.460 ;
        RECT 21.660 -28.090 22.110 -28.040 ;
        RECT 20.020 -28.380 22.110 -28.090 ;
        RECT 20.020 -28.430 20.470 -28.380 ;
        RECT 3.270 -29.010 3.720 -28.940 ;
        RECT 1.420 -29.250 3.720 -29.010 ;
        RECT 1.420 -29.360 1.870 -29.250 ;
        RECT 3.270 -29.360 3.720 -29.250 ;
        RECT 4.670 -29.010 5.120 -28.910 ;
        RECT 6.520 -29.010 6.970 -28.910 ;
        RECT 4.670 -29.250 6.970 -29.010 ;
        RECT 4.670 -29.330 5.120 -29.250 ;
        RECT 5.720 -29.690 6.130 -29.250 ;
        RECT 6.520 -29.360 6.970 -29.250 ;
        RECT 8.160 -29.010 8.610 -28.910 ;
        RECT 10.010 -29.010 10.460 -28.910 ;
        RECT 8.160 -29.250 10.460 -29.010 ;
        RECT 8.160 -29.360 8.610 -29.250 ;
        RECT 9.000 -29.690 9.410 -29.250 ;
        RECT 10.010 -29.330 10.460 -29.250 ;
        RECT 11.410 -29.010 11.860 -28.940 ;
        RECT 12.460 -29.010 12.870 -28.580 ;
        RECT 13.260 -29.010 13.710 -28.910 ;
        RECT 11.410 -29.250 13.710 -29.010 ;
        RECT 11.410 -29.360 11.860 -29.250 ;
        RECT 13.260 -29.360 13.710 -29.250 ;
        RECT 14.920 -29.010 15.370 -28.910 ;
        RECT 15.760 -29.010 16.170 -28.580 ;
        RECT 18.920 -28.650 20.470 -28.430 ;
        RECT 20.850 -28.440 21.280 -28.380 ;
        RECT 21.660 -28.430 22.110 -28.380 ;
        RECT 22.710 -28.430 23.210 -28.040 ;
        RECT 21.660 -28.650 23.210 -28.430 ;
        RECT 32.420 -28.040 33.970 -27.820 ;
        RECT 32.420 -28.430 32.920 -28.040 ;
        RECT 33.520 -28.090 33.970 -28.040 ;
        RECT 34.350 -28.090 34.780 -28.030 ;
        RECT 35.160 -28.040 36.710 -27.820 ;
        RECT 39.460 -27.890 39.870 -27.460 ;
        RECT 40.260 -27.560 40.710 -27.460 ;
        RECT 41.920 -27.220 42.370 -27.110 ;
        RECT 43.770 -27.220 44.220 -27.110 ;
        RECT 41.920 -27.460 44.220 -27.220 ;
        RECT 41.920 -27.560 42.370 -27.460 ;
        RECT 42.760 -27.890 43.170 -27.460 ;
        RECT 43.770 -27.530 44.220 -27.460 ;
        RECT 45.170 -27.220 45.620 -27.140 ;
        RECT 46.220 -27.220 46.630 -26.780 ;
        RECT 47.020 -27.220 47.470 -27.110 ;
        RECT 45.170 -27.460 47.470 -27.220 ;
        RECT 45.170 -27.560 45.620 -27.460 ;
        RECT 47.020 -27.560 47.470 -27.460 ;
        RECT 48.660 -27.220 49.110 -27.110 ;
        RECT 49.500 -27.220 49.910 -26.780 ;
        RECT 52.680 -27.050 53.130 -26.770 ;
        RECT 56.500 -27.050 56.950 -26.770 ;
        RECT 66.180 -26.770 67.710 -26.560 ;
        RECT 68.090 -26.650 68.540 -26.560 ;
        RECT 68.920 -26.770 70.450 -26.560 ;
        RECT 50.510 -27.220 50.960 -27.140 ;
        RECT 48.660 -27.460 50.960 -27.220 ;
        RECT 48.660 -27.560 49.110 -27.460 ;
        RECT 50.510 -27.560 50.960 -27.460 ;
        RECT 51.910 -27.220 52.360 -27.110 ;
        RECT 53.760 -27.220 54.210 -27.110 ;
        RECT 51.910 -27.460 54.210 -27.220 ;
        RECT 51.910 -27.530 52.360 -27.460 ;
        RECT 35.160 -28.090 35.610 -28.040 ;
        RECT 33.520 -28.380 35.610 -28.090 ;
        RECT 33.520 -28.430 33.970 -28.380 ;
        RECT 16.770 -29.010 17.220 -28.940 ;
        RECT 14.920 -29.250 17.220 -29.010 ;
        RECT 14.920 -29.360 15.370 -29.250 ;
        RECT 16.770 -29.360 17.220 -29.250 ;
        RECT 18.170 -29.010 18.620 -28.910 ;
        RECT 20.020 -29.010 20.470 -28.910 ;
        RECT 18.170 -29.250 20.470 -29.010 ;
        RECT 18.170 -29.330 18.620 -29.250 ;
        RECT 12.180 -29.700 12.630 -29.420 ;
        RECT 16.000 -29.700 16.450 -29.420 ;
        RECT 19.220 -29.690 19.630 -29.250 ;
        RECT 20.020 -29.360 20.470 -29.250 ;
        RECT 21.660 -29.010 22.110 -28.910 ;
        RECT 23.510 -29.010 23.960 -28.910 ;
        RECT 21.660 -29.250 23.960 -29.010 ;
        RECT 21.660 -29.360 22.110 -29.250 ;
        RECT 22.500 -29.690 22.910 -29.250 ;
        RECT 23.510 -29.330 23.960 -29.250 ;
        RECT 24.910 -29.010 25.360 -28.940 ;
        RECT 25.960 -29.010 26.370 -28.580 ;
        RECT 26.760 -29.010 27.210 -28.910 ;
        RECT 24.910 -29.250 27.210 -29.010 ;
        RECT 24.910 -29.360 25.360 -29.250 ;
        RECT 26.760 -29.360 27.210 -29.250 ;
        RECT 28.420 -29.010 28.870 -28.910 ;
        RECT 29.260 -29.010 29.670 -28.580 ;
        RECT 32.420 -28.650 33.970 -28.430 ;
        RECT 34.350 -28.440 34.780 -28.380 ;
        RECT 35.160 -28.430 35.610 -28.380 ;
        RECT 36.210 -28.430 36.710 -28.040 ;
        RECT 35.160 -28.650 36.710 -28.430 ;
        RECT 45.920 -28.040 47.470 -27.820 ;
        RECT 45.920 -28.430 46.420 -28.040 ;
        RECT 47.020 -28.090 47.470 -28.040 ;
        RECT 47.850 -28.090 48.280 -28.030 ;
        RECT 48.660 -28.040 50.210 -27.820 ;
        RECT 52.960 -27.890 53.370 -27.460 ;
        RECT 53.760 -27.560 54.210 -27.460 ;
        RECT 55.420 -27.220 55.870 -27.110 ;
        RECT 57.270 -27.220 57.720 -27.110 ;
        RECT 55.420 -27.460 57.720 -27.220 ;
        RECT 55.420 -27.560 55.870 -27.460 ;
        RECT 56.260 -27.890 56.670 -27.460 ;
        RECT 57.270 -27.530 57.720 -27.460 ;
        RECT 58.670 -27.220 59.120 -27.140 ;
        RECT 59.720 -27.220 60.130 -26.780 ;
        RECT 60.520 -27.220 60.970 -27.110 ;
        RECT 58.670 -27.460 60.970 -27.220 ;
        RECT 58.670 -27.560 59.120 -27.460 ;
        RECT 60.520 -27.560 60.970 -27.460 ;
        RECT 62.160 -27.220 62.610 -27.110 ;
        RECT 63.000 -27.220 63.410 -26.780 ;
        RECT 66.180 -27.050 66.630 -26.770 ;
        RECT 70.000 -27.050 70.450 -26.770 ;
        RECT 79.680 -26.770 81.210 -26.560 ;
        RECT 81.590 -26.650 82.040 -26.560 ;
        RECT 82.420 -26.770 83.950 -26.560 ;
        RECT 64.010 -27.220 64.460 -27.140 ;
        RECT 62.160 -27.460 64.460 -27.220 ;
        RECT 62.160 -27.560 62.610 -27.460 ;
        RECT 64.010 -27.560 64.460 -27.460 ;
        RECT 65.410 -27.220 65.860 -27.110 ;
        RECT 67.260 -27.220 67.710 -27.110 ;
        RECT 65.410 -27.460 67.710 -27.220 ;
        RECT 65.410 -27.530 65.860 -27.460 ;
        RECT 48.660 -28.090 49.110 -28.040 ;
        RECT 47.020 -28.380 49.110 -28.090 ;
        RECT 47.020 -28.430 47.470 -28.380 ;
        RECT 30.270 -29.010 30.720 -28.940 ;
        RECT 28.420 -29.250 30.720 -29.010 ;
        RECT 28.420 -29.360 28.870 -29.250 ;
        RECT 30.270 -29.360 30.720 -29.250 ;
        RECT 31.670 -29.010 32.120 -28.910 ;
        RECT 33.520 -29.010 33.970 -28.910 ;
        RECT 31.670 -29.250 33.970 -29.010 ;
        RECT 31.670 -29.330 32.120 -29.250 ;
        RECT 12.180 -29.910 13.710 -29.700 ;
        RECT 14.090 -29.910 14.540 -29.820 ;
        RECT 14.920 -29.910 16.450 -29.700 ;
        RECT 25.680 -29.700 26.130 -29.420 ;
        RECT 29.500 -29.700 29.950 -29.420 ;
        RECT 32.720 -29.690 33.130 -29.250 ;
        RECT 33.520 -29.360 33.970 -29.250 ;
        RECT 35.160 -29.010 35.610 -28.910 ;
        RECT 37.010 -29.010 37.460 -28.910 ;
        RECT 35.160 -29.250 37.460 -29.010 ;
        RECT 35.160 -29.360 35.610 -29.250 ;
        RECT 36.000 -29.690 36.410 -29.250 ;
        RECT 37.010 -29.330 37.460 -29.250 ;
        RECT 38.410 -29.010 38.860 -28.940 ;
        RECT 39.460 -29.010 39.870 -28.580 ;
        RECT 40.260 -29.010 40.710 -28.910 ;
        RECT 38.410 -29.250 40.710 -29.010 ;
        RECT 38.410 -29.360 38.860 -29.250 ;
        RECT 40.260 -29.360 40.710 -29.250 ;
        RECT 41.920 -29.010 42.370 -28.910 ;
        RECT 42.760 -29.010 43.170 -28.580 ;
        RECT 45.920 -28.650 47.470 -28.430 ;
        RECT 47.850 -28.440 48.280 -28.380 ;
        RECT 48.660 -28.430 49.110 -28.380 ;
        RECT 49.710 -28.430 50.210 -28.040 ;
        RECT 48.660 -28.650 50.210 -28.430 ;
        RECT 59.420 -28.040 60.970 -27.820 ;
        RECT 59.420 -28.430 59.920 -28.040 ;
        RECT 60.520 -28.090 60.970 -28.040 ;
        RECT 61.350 -28.090 61.780 -28.030 ;
        RECT 62.160 -28.040 63.710 -27.820 ;
        RECT 66.460 -27.890 66.870 -27.460 ;
        RECT 67.260 -27.560 67.710 -27.460 ;
        RECT 68.920 -27.220 69.370 -27.110 ;
        RECT 70.770 -27.220 71.220 -27.110 ;
        RECT 68.920 -27.460 71.220 -27.220 ;
        RECT 68.920 -27.560 69.370 -27.460 ;
        RECT 69.760 -27.890 70.170 -27.460 ;
        RECT 70.770 -27.530 71.220 -27.460 ;
        RECT 72.170 -27.220 72.620 -27.140 ;
        RECT 73.220 -27.220 73.630 -26.780 ;
        RECT 74.020 -27.220 74.470 -27.110 ;
        RECT 72.170 -27.460 74.470 -27.220 ;
        RECT 72.170 -27.560 72.620 -27.460 ;
        RECT 74.020 -27.560 74.470 -27.460 ;
        RECT 75.660 -27.220 76.110 -27.110 ;
        RECT 76.500 -27.220 76.910 -26.780 ;
        RECT 79.680 -27.050 80.130 -26.770 ;
        RECT 83.500 -27.050 83.950 -26.770 ;
        RECT 93.180 -26.770 94.710 -26.560 ;
        RECT 95.090 -26.650 95.540 -26.560 ;
        RECT 95.920 -26.770 97.450 -26.560 ;
        RECT 77.510 -27.220 77.960 -27.140 ;
        RECT 75.660 -27.460 77.960 -27.220 ;
        RECT 75.660 -27.560 76.110 -27.460 ;
        RECT 77.510 -27.560 77.960 -27.460 ;
        RECT 78.910 -27.220 79.360 -27.110 ;
        RECT 80.760 -27.220 81.210 -27.110 ;
        RECT 78.910 -27.460 81.210 -27.220 ;
        RECT 78.910 -27.530 79.360 -27.460 ;
        RECT 62.160 -28.090 62.610 -28.040 ;
        RECT 60.520 -28.380 62.610 -28.090 ;
        RECT 60.520 -28.430 60.970 -28.380 ;
        RECT 43.770 -29.010 44.220 -28.940 ;
        RECT 41.920 -29.250 44.220 -29.010 ;
        RECT 41.920 -29.360 42.370 -29.250 ;
        RECT 43.770 -29.360 44.220 -29.250 ;
        RECT 45.170 -29.010 45.620 -28.910 ;
        RECT 47.020 -29.010 47.470 -28.910 ;
        RECT 45.170 -29.250 47.470 -29.010 ;
        RECT 45.170 -29.330 45.620 -29.250 ;
        RECT 25.680 -29.910 27.210 -29.700 ;
        RECT 27.590 -29.910 28.040 -29.820 ;
        RECT 28.420 -29.910 29.950 -29.700 ;
        RECT 39.180 -29.700 39.630 -29.420 ;
        RECT 43.000 -29.700 43.450 -29.420 ;
        RECT 46.220 -29.690 46.630 -29.250 ;
        RECT 47.020 -29.360 47.470 -29.250 ;
        RECT 48.660 -29.010 49.110 -28.910 ;
        RECT 50.510 -29.010 50.960 -28.910 ;
        RECT 48.660 -29.250 50.960 -29.010 ;
        RECT 48.660 -29.360 49.110 -29.250 ;
        RECT 49.500 -29.690 49.910 -29.250 ;
        RECT 50.510 -29.330 50.960 -29.250 ;
        RECT 51.910 -29.010 52.360 -28.940 ;
        RECT 52.960 -29.010 53.370 -28.580 ;
        RECT 53.760 -29.010 54.210 -28.910 ;
        RECT 51.910 -29.250 54.210 -29.010 ;
        RECT 51.910 -29.360 52.360 -29.250 ;
        RECT 53.760 -29.360 54.210 -29.250 ;
        RECT 55.420 -29.010 55.870 -28.910 ;
        RECT 56.260 -29.010 56.670 -28.580 ;
        RECT 59.420 -28.650 60.970 -28.430 ;
        RECT 61.350 -28.440 61.780 -28.380 ;
        RECT 62.160 -28.430 62.610 -28.380 ;
        RECT 63.210 -28.430 63.710 -28.040 ;
        RECT 62.160 -28.650 63.710 -28.430 ;
        RECT 72.920 -28.040 74.470 -27.820 ;
        RECT 72.920 -28.430 73.420 -28.040 ;
        RECT 74.020 -28.090 74.470 -28.040 ;
        RECT 74.850 -28.090 75.280 -28.030 ;
        RECT 75.660 -28.040 77.210 -27.820 ;
        RECT 79.960 -27.890 80.370 -27.460 ;
        RECT 80.760 -27.560 81.210 -27.460 ;
        RECT 82.420 -27.220 82.870 -27.110 ;
        RECT 84.270 -27.220 84.720 -27.110 ;
        RECT 82.420 -27.460 84.720 -27.220 ;
        RECT 82.420 -27.560 82.870 -27.460 ;
        RECT 83.260 -27.890 83.670 -27.460 ;
        RECT 84.270 -27.530 84.720 -27.460 ;
        RECT 85.670 -27.220 86.120 -27.140 ;
        RECT 86.720 -27.220 87.130 -26.780 ;
        RECT 87.520 -27.220 87.970 -27.110 ;
        RECT 85.670 -27.460 87.970 -27.220 ;
        RECT 85.670 -27.560 86.120 -27.460 ;
        RECT 87.520 -27.560 87.970 -27.460 ;
        RECT 89.160 -27.220 89.610 -27.110 ;
        RECT 90.000 -27.220 90.410 -26.780 ;
        RECT 93.180 -27.050 93.630 -26.770 ;
        RECT 97.000 -27.050 97.450 -26.770 ;
        RECT 106.680 -26.610 110.950 -26.560 ;
        RECT 106.680 -26.770 108.210 -26.610 ;
        RECT 108.590 -26.650 109.040 -26.610 ;
        RECT 109.420 -26.770 110.950 -26.610 ;
        RECT 91.010 -27.220 91.460 -27.140 ;
        RECT 89.160 -27.460 91.460 -27.220 ;
        RECT 89.160 -27.560 89.610 -27.460 ;
        RECT 91.010 -27.560 91.460 -27.460 ;
        RECT 92.410 -27.220 92.860 -27.110 ;
        RECT 94.260 -27.220 94.710 -27.110 ;
        RECT 92.410 -27.460 94.710 -27.220 ;
        RECT 92.410 -27.530 92.860 -27.460 ;
        RECT 75.660 -28.090 76.110 -28.040 ;
        RECT 74.020 -28.380 76.110 -28.090 ;
        RECT 74.020 -28.430 74.470 -28.380 ;
        RECT 57.270 -29.010 57.720 -28.940 ;
        RECT 55.420 -29.250 57.720 -29.010 ;
        RECT 55.420 -29.360 55.870 -29.250 ;
        RECT 57.270 -29.360 57.720 -29.250 ;
        RECT 58.670 -29.010 59.120 -28.910 ;
        RECT 60.520 -29.010 60.970 -28.910 ;
        RECT 58.670 -29.250 60.970 -29.010 ;
        RECT 58.670 -29.330 59.120 -29.250 ;
        RECT 39.180 -29.910 40.710 -29.700 ;
        RECT 41.090 -29.910 41.540 -29.820 ;
        RECT 41.920 -29.910 43.450 -29.700 ;
        RECT 52.680 -29.700 53.130 -29.420 ;
        RECT 56.500 -29.700 56.950 -29.420 ;
        RECT 59.720 -29.690 60.130 -29.250 ;
        RECT 60.520 -29.360 60.970 -29.250 ;
        RECT 62.160 -29.010 62.610 -28.910 ;
        RECT 64.010 -29.010 64.460 -28.910 ;
        RECT 62.160 -29.250 64.460 -29.010 ;
        RECT 62.160 -29.360 62.610 -29.250 ;
        RECT 63.000 -29.690 63.410 -29.250 ;
        RECT 64.010 -29.330 64.460 -29.250 ;
        RECT 65.410 -29.010 65.860 -28.940 ;
        RECT 66.460 -29.010 66.870 -28.580 ;
        RECT 67.260 -29.010 67.710 -28.910 ;
        RECT 65.410 -29.250 67.710 -29.010 ;
        RECT 65.410 -29.360 65.860 -29.250 ;
        RECT 67.260 -29.360 67.710 -29.250 ;
        RECT 68.920 -29.010 69.370 -28.910 ;
        RECT 69.760 -29.010 70.170 -28.580 ;
        RECT 72.920 -28.650 74.470 -28.430 ;
        RECT 74.850 -28.440 75.280 -28.380 ;
        RECT 75.660 -28.430 76.110 -28.380 ;
        RECT 76.710 -28.430 77.210 -28.040 ;
        RECT 75.660 -28.650 77.210 -28.430 ;
        RECT 86.420 -28.040 87.970 -27.820 ;
        RECT 86.420 -28.430 86.920 -28.040 ;
        RECT 87.520 -28.090 87.970 -28.040 ;
        RECT 88.350 -28.090 88.780 -28.030 ;
        RECT 89.160 -28.040 90.710 -27.820 ;
        RECT 93.460 -27.890 93.870 -27.460 ;
        RECT 94.260 -27.560 94.710 -27.460 ;
        RECT 95.920 -27.220 96.370 -27.110 ;
        RECT 97.770 -27.220 98.220 -27.110 ;
        RECT 95.920 -27.460 98.220 -27.220 ;
        RECT 95.920 -27.560 96.370 -27.460 ;
        RECT 96.760 -27.890 97.170 -27.460 ;
        RECT 97.770 -27.530 98.220 -27.460 ;
        RECT 99.170 -27.220 99.620 -27.140 ;
        RECT 100.220 -27.220 100.630 -26.780 ;
        RECT 101.020 -27.220 101.470 -27.110 ;
        RECT 99.170 -27.460 101.470 -27.220 ;
        RECT 99.170 -27.560 99.620 -27.460 ;
        RECT 101.020 -27.560 101.470 -27.460 ;
        RECT 102.660 -27.220 103.110 -27.110 ;
        RECT 103.500 -27.220 103.910 -26.780 ;
        RECT 106.680 -27.050 107.130 -26.770 ;
        RECT 110.500 -27.050 110.950 -26.770 ;
        RECT 120.180 -26.770 121.710 -26.560 ;
        RECT 122.090 -26.650 122.540 -26.560 ;
        RECT 122.920 -26.770 124.450 -26.560 ;
        RECT 104.510 -27.220 104.960 -27.140 ;
        RECT 102.660 -27.460 104.960 -27.220 ;
        RECT 102.660 -27.560 103.110 -27.460 ;
        RECT 104.510 -27.560 104.960 -27.460 ;
        RECT 105.910 -27.220 106.360 -27.110 ;
        RECT 107.760 -27.220 108.210 -27.110 ;
        RECT 105.910 -27.460 108.210 -27.220 ;
        RECT 105.910 -27.530 106.360 -27.460 ;
        RECT 89.160 -28.090 89.610 -28.040 ;
        RECT 87.520 -28.380 89.610 -28.090 ;
        RECT 87.520 -28.430 87.970 -28.380 ;
        RECT 70.770 -29.010 71.220 -28.940 ;
        RECT 68.920 -29.250 71.220 -29.010 ;
        RECT 68.920 -29.360 69.370 -29.250 ;
        RECT 70.770 -29.360 71.220 -29.250 ;
        RECT 72.170 -29.010 72.620 -28.910 ;
        RECT 74.020 -29.010 74.470 -28.910 ;
        RECT 72.170 -29.250 74.470 -29.010 ;
        RECT 72.170 -29.330 72.620 -29.250 ;
        RECT 52.680 -29.910 54.210 -29.700 ;
        RECT 54.590 -29.910 55.040 -29.820 ;
        RECT 55.420 -29.910 56.950 -29.700 ;
        RECT 66.180 -29.700 66.630 -29.420 ;
        RECT 70.000 -29.700 70.450 -29.420 ;
        RECT 73.220 -29.690 73.630 -29.250 ;
        RECT 74.020 -29.360 74.470 -29.250 ;
        RECT 75.660 -29.010 76.110 -28.910 ;
        RECT 77.510 -29.010 77.960 -28.910 ;
        RECT 75.660 -29.250 77.960 -29.010 ;
        RECT 75.660 -29.360 76.110 -29.250 ;
        RECT 76.500 -29.690 76.910 -29.250 ;
        RECT 77.510 -29.330 77.960 -29.250 ;
        RECT 78.910 -29.010 79.360 -28.940 ;
        RECT 79.960 -29.010 80.370 -28.580 ;
        RECT 80.760 -29.010 81.210 -28.910 ;
        RECT 78.910 -29.250 81.210 -29.010 ;
        RECT 78.910 -29.360 79.360 -29.250 ;
        RECT 80.760 -29.360 81.210 -29.250 ;
        RECT 82.420 -29.010 82.870 -28.910 ;
        RECT 83.260 -29.010 83.670 -28.580 ;
        RECT 86.420 -28.650 87.970 -28.430 ;
        RECT 88.350 -28.440 88.780 -28.380 ;
        RECT 89.160 -28.430 89.610 -28.380 ;
        RECT 90.210 -28.430 90.710 -28.040 ;
        RECT 89.160 -28.650 90.710 -28.430 ;
        RECT 99.920 -28.040 101.470 -27.820 ;
        RECT 99.920 -28.430 100.420 -28.040 ;
        RECT 101.020 -28.090 101.470 -28.040 ;
        RECT 101.850 -28.090 102.280 -28.030 ;
        RECT 102.660 -28.040 104.210 -27.820 ;
        RECT 106.960 -27.890 107.370 -27.460 ;
        RECT 107.760 -27.560 108.210 -27.460 ;
        RECT 109.420 -27.220 109.870 -27.110 ;
        RECT 111.270 -27.220 111.720 -27.110 ;
        RECT 109.420 -27.460 111.720 -27.220 ;
        RECT 109.420 -27.560 109.870 -27.460 ;
        RECT 110.260 -27.890 110.670 -27.460 ;
        RECT 111.270 -27.530 111.720 -27.460 ;
        RECT 112.670 -27.220 113.120 -27.140 ;
        RECT 113.720 -27.220 114.130 -26.780 ;
        RECT 114.520 -27.220 114.970 -27.110 ;
        RECT 112.670 -27.460 114.970 -27.220 ;
        RECT 112.670 -27.560 113.120 -27.460 ;
        RECT 114.520 -27.560 114.970 -27.460 ;
        RECT 116.160 -27.220 116.610 -27.110 ;
        RECT 117.000 -27.220 117.410 -26.780 ;
        RECT 120.180 -27.050 120.630 -26.770 ;
        RECT 124.000 -27.050 124.450 -26.770 ;
        RECT 133.680 -26.770 135.210 -26.560 ;
        RECT 135.590 -26.650 136.040 -26.560 ;
        RECT 136.420 -26.770 137.950 -26.560 ;
        RECT 118.010 -27.220 118.460 -27.140 ;
        RECT 116.160 -27.460 118.460 -27.220 ;
        RECT 116.160 -27.560 116.610 -27.460 ;
        RECT 118.010 -27.560 118.460 -27.460 ;
        RECT 119.410 -27.220 119.860 -27.110 ;
        RECT 121.260 -27.220 121.710 -27.110 ;
        RECT 119.410 -27.460 121.710 -27.220 ;
        RECT 119.410 -27.530 119.860 -27.460 ;
        RECT 102.660 -28.090 103.110 -28.040 ;
        RECT 101.020 -28.380 103.110 -28.090 ;
        RECT 101.020 -28.430 101.470 -28.380 ;
        RECT 84.270 -29.010 84.720 -28.940 ;
        RECT 82.420 -29.250 84.720 -29.010 ;
        RECT 82.420 -29.360 82.870 -29.250 ;
        RECT 84.270 -29.360 84.720 -29.250 ;
        RECT 85.670 -29.010 86.120 -28.910 ;
        RECT 87.520 -29.010 87.970 -28.910 ;
        RECT 85.670 -29.250 87.970 -29.010 ;
        RECT 85.670 -29.330 86.120 -29.250 ;
        RECT 66.180 -29.910 67.710 -29.700 ;
        RECT 68.090 -29.910 68.540 -29.820 ;
        RECT 68.920 -29.910 70.450 -29.700 ;
        RECT 79.680 -29.700 80.130 -29.420 ;
        RECT 83.500 -29.700 83.950 -29.420 ;
        RECT 86.720 -29.690 87.130 -29.250 ;
        RECT 87.520 -29.360 87.970 -29.250 ;
        RECT 89.160 -29.010 89.610 -28.910 ;
        RECT 91.010 -29.010 91.460 -28.910 ;
        RECT 89.160 -29.250 91.460 -29.010 ;
        RECT 89.160 -29.360 89.610 -29.250 ;
        RECT 90.000 -29.690 90.410 -29.250 ;
        RECT 91.010 -29.330 91.460 -29.250 ;
        RECT 92.410 -29.010 92.860 -28.940 ;
        RECT 93.460 -29.010 93.870 -28.580 ;
        RECT 94.260 -29.010 94.710 -28.910 ;
        RECT 92.410 -29.250 94.710 -29.010 ;
        RECT 92.410 -29.360 92.860 -29.250 ;
        RECT 94.260 -29.360 94.710 -29.250 ;
        RECT 95.920 -29.010 96.370 -28.910 ;
        RECT 96.760 -29.010 97.170 -28.580 ;
        RECT 99.920 -28.650 101.470 -28.430 ;
        RECT 101.850 -28.440 102.280 -28.380 ;
        RECT 102.660 -28.430 103.110 -28.380 ;
        RECT 103.710 -28.430 104.210 -28.040 ;
        RECT 102.660 -28.650 104.210 -28.430 ;
        RECT 113.420 -28.040 114.970 -27.820 ;
        RECT 113.420 -28.430 113.920 -28.040 ;
        RECT 114.520 -28.090 114.970 -28.040 ;
        RECT 115.350 -28.090 115.780 -28.030 ;
        RECT 116.160 -28.040 117.710 -27.820 ;
        RECT 120.460 -27.890 120.870 -27.460 ;
        RECT 121.260 -27.560 121.710 -27.460 ;
        RECT 122.920 -27.220 123.370 -27.110 ;
        RECT 124.770 -27.220 125.220 -27.110 ;
        RECT 122.920 -27.460 125.220 -27.220 ;
        RECT 122.920 -27.560 123.370 -27.460 ;
        RECT 123.760 -27.890 124.170 -27.460 ;
        RECT 124.770 -27.530 125.220 -27.460 ;
        RECT 126.170 -27.220 126.620 -27.140 ;
        RECT 127.220 -27.220 127.630 -26.780 ;
        RECT 128.020 -27.220 128.470 -27.110 ;
        RECT 126.170 -27.460 128.470 -27.220 ;
        RECT 126.170 -27.560 126.620 -27.460 ;
        RECT 128.020 -27.560 128.470 -27.460 ;
        RECT 129.660 -27.220 130.110 -27.110 ;
        RECT 130.500 -27.220 130.910 -26.780 ;
        RECT 133.680 -27.050 134.130 -26.770 ;
        RECT 137.500 -27.050 137.950 -26.770 ;
        RECT 147.180 -26.770 148.710 -26.560 ;
        RECT 149.090 -26.650 149.540 -26.560 ;
        RECT 149.920 -26.770 151.450 -26.560 ;
        RECT 131.510 -27.220 131.960 -27.140 ;
        RECT 129.660 -27.460 131.960 -27.220 ;
        RECT 129.660 -27.560 130.110 -27.460 ;
        RECT 131.510 -27.560 131.960 -27.460 ;
        RECT 132.910 -27.220 133.360 -27.110 ;
        RECT 134.760 -27.220 135.210 -27.110 ;
        RECT 132.910 -27.460 135.210 -27.220 ;
        RECT 132.910 -27.530 133.360 -27.460 ;
        RECT 116.160 -28.090 116.610 -28.040 ;
        RECT 114.520 -28.380 116.610 -28.090 ;
        RECT 114.520 -28.430 114.970 -28.380 ;
        RECT 97.770 -29.010 98.220 -28.940 ;
        RECT 95.920 -29.250 98.220 -29.010 ;
        RECT 95.920 -29.360 96.370 -29.250 ;
        RECT 97.770 -29.360 98.220 -29.250 ;
        RECT 99.170 -29.010 99.620 -28.910 ;
        RECT 101.020 -29.010 101.470 -28.910 ;
        RECT 99.170 -29.250 101.470 -29.010 ;
        RECT 99.170 -29.330 99.620 -29.250 ;
        RECT 79.680 -29.910 81.210 -29.700 ;
        RECT 81.590 -29.910 82.040 -29.820 ;
        RECT 82.420 -29.910 83.950 -29.700 ;
        RECT 93.180 -29.700 93.630 -29.420 ;
        RECT 97.000 -29.700 97.450 -29.420 ;
        RECT 100.220 -29.690 100.630 -29.250 ;
        RECT 101.020 -29.360 101.470 -29.250 ;
        RECT 102.660 -29.010 103.110 -28.910 ;
        RECT 104.510 -29.010 104.960 -28.910 ;
        RECT 102.660 -29.250 104.960 -29.010 ;
        RECT 102.660 -29.360 103.110 -29.250 ;
        RECT 103.500 -29.690 103.910 -29.250 ;
        RECT 104.510 -29.330 104.960 -29.250 ;
        RECT 105.910 -29.010 106.360 -28.940 ;
        RECT 106.960 -29.010 107.370 -28.580 ;
        RECT 107.760 -29.010 108.210 -28.910 ;
        RECT 105.910 -29.250 108.210 -29.010 ;
        RECT 105.910 -29.360 106.360 -29.250 ;
        RECT 107.760 -29.360 108.210 -29.250 ;
        RECT 109.420 -29.010 109.870 -28.910 ;
        RECT 110.260 -29.010 110.670 -28.580 ;
        RECT 113.420 -28.650 114.970 -28.430 ;
        RECT 115.350 -28.440 115.780 -28.380 ;
        RECT 116.160 -28.430 116.610 -28.380 ;
        RECT 117.210 -28.430 117.710 -28.040 ;
        RECT 116.160 -28.650 117.710 -28.430 ;
        RECT 126.920 -28.040 128.470 -27.820 ;
        RECT 126.920 -28.430 127.420 -28.040 ;
        RECT 128.020 -28.090 128.470 -28.040 ;
        RECT 128.850 -28.090 129.280 -28.030 ;
        RECT 129.660 -28.040 131.210 -27.820 ;
        RECT 133.960 -27.890 134.370 -27.460 ;
        RECT 134.760 -27.560 135.210 -27.460 ;
        RECT 136.420 -27.220 136.870 -27.110 ;
        RECT 138.270 -27.220 138.720 -27.110 ;
        RECT 136.420 -27.460 138.720 -27.220 ;
        RECT 136.420 -27.560 136.870 -27.460 ;
        RECT 137.260 -27.890 137.670 -27.460 ;
        RECT 138.270 -27.530 138.720 -27.460 ;
        RECT 139.670 -27.220 140.120 -27.140 ;
        RECT 140.720 -27.220 141.130 -26.780 ;
        RECT 141.520 -27.220 141.970 -27.110 ;
        RECT 139.670 -27.460 141.970 -27.220 ;
        RECT 139.670 -27.560 140.120 -27.460 ;
        RECT 141.520 -27.560 141.970 -27.460 ;
        RECT 143.160 -27.220 143.610 -27.110 ;
        RECT 144.000 -27.220 144.410 -26.780 ;
        RECT 147.180 -27.050 147.630 -26.770 ;
        RECT 151.000 -27.050 151.450 -26.770 ;
        RECT 160.680 -26.610 164.950 -26.560 ;
        RECT 160.680 -26.770 162.210 -26.610 ;
        RECT 162.590 -26.650 163.040 -26.610 ;
        RECT 163.420 -26.770 164.950 -26.610 ;
        RECT 145.010 -27.220 145.460 -27.140 ;
        RECT 143.160 -27.460 145.460 -27.220 ;
        RECT 143.160 -27.560 143.610 -27.460 ;
        RECT 145.010 -27.560 145.460 -27.460 ;
        RECT 146.410 -27.220 146.860 -27.110 ;
        RECT 148.260 -27.220 148.710 -27.110 ;
        RECT 146.410 -27.460 148.710 -27.220 ;
        RECT 146.410 -27.530 146.860 -27.460 ;
        RECT 129.660 -28.090 130.110 -28.040 ;
        RECT 128.020 -28.380 130.110 -28.090 ;
        RECT 128.020 -28.430 128.470 -28.380 ;
        RECT 111.270 -29.010 111.720 -28.940 ;
        RECT 109.420 -29.250 111.720 -29.010 ;
        RECT 109.420 -29.360 109.870 -29.250 ;
        RECT 111.270 -29.360 111.720 -29.250 ;
        RECT 112.670 -29.010 113.120 -28.910 ;
        RECT 114.520 -29.010 114.970 -28.910 ;
        RECT 112.670 -29.250 114.970 -29.010 ;
        RECT 112.670 -29.330 113.120 -29.250 ;
        RECT 93.180 -29.910 94.710 -29.700 ;
        RECT 95.090 -29.910 95.540 -29.820 ;
        RECT 95.920 -29.910 97.450 -29.700 ;
        RECT 106.680 -29.700 107.130 -29.420 ;
        RECT 110.500 -29.700 110.950 -29.420 ;
        RECT 113.720 -29.690 114.130 -29.250 ;
        RECT 114.520 -29.360 114.970 -29.250 ;
        RECT 116.160 -29.010 116.610 -28.910 ;
        RECT 118.010 -29.010 118.460 -28.910 ;
        RECT 116.160 -29.250 118.460 -29.010 ;
        RECT 116.160 -29.360 116.610 -29.250 ;
        RECT 117.000 -29.690 117.410 -29.250 ;
        RECT 118.010 -29.330 118.460 -29.250 ;
        RECT 119.410 -29.010 119.860 -28.940 ;
        RECT 120.460 -29.010 120.870 -28.580 ;
        RECT 121.260 -29.010 121.710 -28.910 ;
        RECT 119.410 -29.250 121.710 -29.010 ;
        RECT 119.410 -29.360 119.860 -29.250 ;
        RECT 121.260 -29.360 121.710 -29.250 ;
        RECT 122.920 -29.010 123.370 -28.910 ;
        RECT 123.760 -29.010 124.170 -28.580 ;
        RECT 126.920 -28.650 128.470 -28.430 ;
        RECT 128.850 -28.440 129.280 -28.380 ;
        RECT 129.660 -28.430 130.110 -28.380 ;
        RECT 130.710 -28.430 131.210 -28.040 ;
        RECT 129.660 -28.650 131.210 -28.430 ;
        RECT 140.420 -28.040 141.970 -27.820 ;
        RECT 140.420 -28.430 140.920 -28.040 ;
        RECT 141.520 -28.090 141.970 -28.040 ;
        RECT 142.350 -28.090 142.780 -28.030 ;
        RECT 143.160 -28.040 144.710 -27.820 ;
        RECT 147.460 -27.890 147.870 -27.460 ;
        RECT 148.260 -27.560 148.710 -27.460 ;
        RECT 149.920 -27.220 150.370 -27.110 ;
        RECT 151.770 -27.220 152.220 -27.110 ;
        RECT 149.920 -27.460 152.220 -27.220 ;
        RECT 149.920 -27.560 150.370 -27.460 ;
        RECT 150.760 -27.890 151.170 -27.460 ;
        RECT 151.770 -27.530 152.220 -27.460 ;
        RECT 153.170 -27.220 153.620 -27.140 ;
        RECT 154.220 -27.220 154.630 -26.780 ;
        RECT 155.020 -27.220 155.470 -27.110 ;
        RECT 153.170 -27.460 155.470 -27.220 ;
        RECT 153.170 -27.560 153.620 -27.460 ;
        RECT 155.020 -27.560 155.470 -27.460 ;
        RECT 156.660 -27.220 157.110 -27.110 ;
        RECT 157.500 -27.220 157.910 -26.780 ;
        RECT 160.680 -27.050 161.130 -26.770 ;
        RECT 164.500 -27.050 164.950 -26.770 ;
        RECT 174.180 -26.770 175.710 -26.560 ;
        RECT 176.090 -26.650 176.540 -26.560 ;
        RECT 176.920 -26.770 178.450 -26.560 ;
        RECT 158.510 -27.220 158.960 -27.140 ;
        RECT 156.660 -27.460 158.960 -27.220 ;
        RECT 156.660 -27.560 157.110 -27.460 ;
        RECT 158.510 -27.560 158.960 -27.460 ;
        RECT 159.910 -27.220 160.360 -27.110 ;
        RECT 161.760 -27.220 162.210 -27.110 ;
        RECT 159.910 -27.460 162.210 -27.220 ;
        RECT 159.910 -27.530 160.360 -27.460 ;
        RECT 143.160 -28.090 143.610 -28.040 ;
        RECT 141.520 -28.380 143.610 -28.090 ;
        RECT 141.520 -28.430 141.970 -28.380 ;
        RECT 124.770 -29.010 125.220 -28.940 ;
        RECT 122.920 -29.250 125.220 -29.010 ;
        RECT 122.920 -29.360 123.370 -29.250 ;
        RECT 124.770 -29.360 125.220 -29.250 ;
        RECT 126.170 -29.010 126.620 -28.910 ;
        RECT 128.020 -29.010 128.470 -28.910 ;
        RECT 126.170 -29.250 128.470 -29.010 ;
        RECT 126.170 -29.330 126.620 -29.250 ;
        RECT 106.680 -29.910 108.210 -29.700 ;
        RECT 108.590 -29.910 109.040 -29.820 ;
        RECT 109.420 -29.910 110.950 -29.700 ;
        RECT 120.180 -29.700 120.630 -29.420 ;
        RECT 124.000 -29.700 124.450 -29.420 ;
        RECT 127.220 -29.690 127.630 -29.250 ;
        RECT 128.020 -29.360 128.470 -29.250 ;
        RECT 129.660 -29.010 130.110 -28.910 ;
        RECT 131.510 -29.010 131.960 -28.910 ;
        RECT 129.660 -29.250 131.960 -29.010 ;
        RECT 129.660 -29.360 130.110 -29.250 ;
        RECT 130.500 -29.690 130.910 -29.250 ;
        RECT 131.510 -29.330 131.960 -29.250 ;
        RECT 132.910 -29.010 133.360 -28.940 ;
        RECT 133.960 -29.010 134.370 -28.580 ;
        RECT 134.760 -29.010 135.210 -28.910 ;
        RECT 132.910 -29.250 135.210 -29.010 ;
        RECT 132.910 -29.360 133.360 -29.250 ;
        RECT 134.760 -29.360 135.210 -29.250 ;
        RECT 136.420 -29.010 136.870 -28.910 ;
        RECT 137.260 -29.010 137.670 -28.580 ;
        RECT 140.420 -28.650 141.970 -28.430 ;
        RECT 142.350 -28.440 142.780 -28.380 ;
        RECT 143.160 -28.430 143.610 -28.380 ;
        RECT 144.210 -28.430 144.710 -28.040 ;
        RECT 143.160 -28.650 144.710 -28.430 ;
        RECT 153.920 -28.040 155.470 -27.820 ;
        RECT 153.920 -28.430 154.420 -28.040 ;
        RECT 155.020 -28.090 155.470 -28.040 ;
        RECT 155.850 -28.090 156.280 -28.030 ;
        RECT 156.660 -28.040 158.210 -27.820 ;
        RECT 160.960 -27.890 161.370 -27.460 ;
        RECT 161.760 -27.560 162.210 -27.460 ;
        RECT 163.420 -27.220 163.870 -27.110 ;
        RECT 165.270 -27.220 165.720 -27.110 ;
        RECT 163.420 -27.460 165.720 -27.220 ;
        RECT 163.420 -27.560 163.870 -27.460 ;
        RECT 164.260 -27.890 164.670 -27.460 ;
        RECT 165.270 -27.530 165.720 -27.460 ;
        RECT 166.670 -27.220 167.120 -27.140 ;
        RECT 167.720 -27.220 168.130 -26.780 ;
        RECT 168.520 -27.220 168.970 -27.110 ;
        RECT 166.670 -27.460 168.970 -27.220 ;
        RECT 166.670 -27.560 167.120 -27.460 ;
        RECT 168.520 -27.560 168.970 -27.460 ;
        RECT 170.160 -27.220 170.610 -27.110 ;
        RECT 171.000 -27.220 171.410 -26.780 ;
        RECT 174.180 -27.050 174.630 -26.770 ;
        RECT 178.000 -27.050 178.450 -26.770 ;
        RECT 187.680 -26.770 189.210 -26.560 ;
        RECT 189.590 -26.650 190.040 -26.560 ;
        RECT 190.420 -26.770 191.950 -26.560 ;
        RECT 172.010 -27.220 172.460 -27.140 ;
        RECT 170.160 -27.460 172.460 -27.220 ;
        RECT 170.160 -27.560 170.610 -27.460 ;
        RECT 172.010 -27.560 172.460 -27.460 ;
        RECT 173.410 -27.220 173.860 -27.110 ;
        RECT 175.260 -27.220 175.710 -27.110 ;
        RECT 173.410 -27.460 175.710 -27.220 ;
        RECT 173.410 -27.530 173.860 -27.460 ;
        RECT 156.660 -28.090 157.110 -28.040 ;
        RECT 155.020 -28.380 157.110 -28.090 ;
        RECT 155.020 -28.430 155.470 -28.380 ;
        RECT 138.270 -29.010 138.720 -28.940 ;
        RECT 136.420 -29.250 138.720 -29.010 ;
        RECT 136.420 -29.360 136.870 -29.250 ;
        RECT 138.270 -29.360 138.720 -29.250 ;
        RECT 139.670 -29.010 140.120 -28.910 ;
        RECT 141.520 -29.010 141.970 -28.910 ;
        RECT 139.670 -29.250 141.970 -29.010 ;
        RECT 139.670 -29.330 140.120 -29.250 ;
        RECT 120.180 -29.910 121.710 -29.700 ;
        RECT 122.090 -29.910 122.540 -29.820 ;
        RECT 122.920 -29.910 124.450 -29.700 ;
        RECT 133.680 -29.700 134.130 -29.420 ;
        RECT 137.500 -29.700 137.950 -29.420 ;
        RECT 140.720 -29.690 141.130 -29.250 ;
        RECT 141.520 -29.360 141.970 -29.250 ;
        RECT 143.160 -29.010 143.610 -28.910 ;
        RECT 145.010 -29.010 145.460 -28.910 ;
        RECT 143.160 -29.250 145.460 -29.010 ;
        RECT 143.160 -29.360 143.610 -29.250 ;
        RECT 144.000 -29.690 144.410 -29.250 ;
        RECT 145.010 -29.330 145.460 -29.250 ;
        RECT 146.410 -29.010 146.860 -28.940 ;
        RECT 147.460 -29.010 147.870 -28.580 ;
        RECT 148.260 -29.010 148.710 -28.910 ;
        RECT 146.410 -29.250 148.710 -29.010 ;
        RECT 146.410 -29.360 146.860 -29.250 ;
        RECT 148.260 -29.360 148.710 -29.250 ;
        RECT 149.920 -29.010 150.370 -28.910 ;
        RECT 150.760 -29.010 151.170 -28.580 ;
        RECT 153.920 -28.650 155.470 -28.430 ;
        RECT 155.850 -28.440 156.280 -28.380 ;
        RECT 156.660 -28.430 157.110 -28.380 ;
        RECT 157.710 -28.430 158.210 -28.040 ;
        RECT 156.660 -28.650 158.210 -28.430 ;
        RECT 167.420 -28.040 168.970 -27.820 ;
        RECT 167.420 -28.430 167.920 -28.040 ;
        RECT 168.520 -28.090 168.970 -28.040 ;
        RECT 169.350 -28.090 169.780 -28.030 ;
        RECT 170.160 -28.040 171.710 -27.820 ;
        RECT 174.460 -27.890 174.870 -27.460 ;
        RECT 175.260 -27.560 175.710 -27.460 ;
        RECT 176.920 -27.220 177.370 -27.110 ;
        RECT 178.770 -27.220 179.220 -27.110 ;
        RECT 176.920 -27.460 179.220 -27.220 ;
        RECT 176.920 -27.560 177.370 -27.460 ;
        RECT 177.760 -27.890 178.170 -27.460 ;
        RECT 178.770 -27.530 179.220 -27.460 ;
        RECT 180.170 -27.220 180.620 -27.140 ;
        RECT 181.220 -27.220 181.630 -26.780 ;
        RECT 182.020 -27.220 182.470 -27.110 ;
        RECT 180.170 -27.460 182.470 -27.220 ;
        RECT 180.170 -27.560 180.620 -27.460 ;
        RECT 182.020 -27.560 182.470 -27.460 ;
        RECT 183.660 -27.220 184.110 -27.110 ;
        RECT 184.500 -27.220 184.910 -26.780 ;
        RECT 187.680 -27.050 188.130 -26.770 ;
        RECT 191.500 -27.050 191.950 -26.770 ;
        RECT 201.180 -26.770 202.710 -26.560 ;
        RECT 203.090 -26.650 203.540 -26.560 ;
        RECT 203.920 -26.770 205.450 -26.560 ;
        RECT 185.510 -27.220 185.960 -27.140 ;
        RECT 183.660 -27.460 185.960 -27.220 ;
        RECT 183.660 -27.560 184.110 -27.460 ;
        RECT 185.510 -27.560 185.960 -27.460 ;
        RECT 186.910 -27.220 187.360 -27.110 ;
        RECT 188.760 -27.220 189.210 -27.110 ;
        RECT 186.910 -27.460 189.210 -27.220 ;
        RECT 186.910 -27.530 187.360 -27.460 ;
        RECT 170.160 -28.090 170.610 -28.040 ;
        RECT 168.520 -28.380 170.610 -28.090 ;
        RECT 168.520 -28.430 168.970 -28.380 ;
        RECT 151.770 -29.010 152.220 -28.940 ;
        RECT 149.920 -29.250 152.220 -29.010 ;
        RECT 149.920 -29.360 150.370 -29.250 ;
        RECT 151.770 -29.360 152.220 -29.250 ;
        RECT 153.170 -29.010 153.620 -28.910 ;
        RECT 155.020 -29.010 155.470 -28.910 ;
        RECT 153.170 -29.250 155.470 -29.010 ;
        RECT 153.170 -29.330 153.620 -29.250 ;
        RECT 133.680 -29.910 135.210 -29.700 ;
        RECT 135.590 -29.910 136.040 -29.820 ;
        RECT 136.420 -29.910 137.950 -29.700 ;
        RECT 147.180 -29.700 147.630 -29.420 ;
        RECT 151.000 -29.700 151.450 -29.420 ;
        RECT 154.220 -29.690 154.630 -29.250 ;
        RECT 155.020 -29.360 155.470 -29.250 ;
        RECT 156.660 -29.010 157.110 -28.910 ;
        RECT 158.510 -29.010 158.960 -28.910 ;
        RECT 156.660 -29.250 158.960 -29.010 ;
        RECT 156.660 -29.360 157.110 -29.250 ;
        RECT 157.500 -29.690 157.910 -29.250 ;
        RECT 158.510 -29.330 158.960 -29.250 ;
        RECT 159.910 -29.010 160.360 -28.940 ;
        RECT 160.960 -29.010 161.370 -28.580 ;
        RECT 161.760 -29.010 162.210 -28.910 ;
        RECT 159.910 -29.250 162.210 -29.010 ;
        RECT 159.910 -29.360 160.360 -29.250 ;
        RECT 161.760 -29.360 162.210 -29.250 ;
        RECT 163.420 -29.010 163.870 -28.910 ;
        RECT 164.260 -29.010 164.670 -28.580 ;
        RECT 167.420 -28.650 168.970 -28.430 ;
        RECT 169.350 -28.440 169.780 -28.380 ;
        RECT 170.160 -28.430 170.610 -28.380 ;
        RECT 171.210 -28.430 171.710 -28.040 ;
        RECT 170.160 -28.650 171.710 -28.430 ;
        RECT 180.920 -28.040 182.470 -27.820 ;
        RECT 180.920 -28.430 181.420 -28.040 ;
        RECT 182.020 -28.090 182.470 -28.040 ;
        RECT 182.850 -28.090 183.280 -28.030 ;
        RECT 183.660 -28.040 185.210 -27.820 ;
        RECT 187.960 -27.890 188.370 -27.460 ;
        RECT 188.760 -27.560 189.210 -27.460 ;
        RECT 190.420 -27.220 190.870 -27.110 ;
        RECT 192.270 -27.220 192.720 -27.110 ;
        RECT 190.420 -27.460 192.720 -27.220 ;
        RECT 190.420 -27.560 190.870 -27.460 ;
        RECT 191.260 -27.890 191.670 -27.460 ;
        RECT 192.270 -27.530 192.720 -27.460 ;
        RECT 193.670 -27.220 194.120 -27.140 ;
        RECT 194.720 -27.220 195.130 -26.780 ;
        RECT 195.520 -27.220 195.970 -27.110 ;
        RECT 193.670 -27.460 195.970 -27.220 ;
        RECT 193.670 -27.560 194.120 -27.460 ;
        RECT 195.520 -27.560 195.970 -27.460 ;
        RECT 197.160 -27.220 197.610 -27.110 ;
        RECT 198.000 -27.220 198.410 -26.780 ;
        RECT 201.180 -27.050 201.630 -26.770 ;
        RECT 205.000 -27.050 205.450 -26.770 ;
        RECT 214.680 -26.770 216.210 -26.560 ;
        RECT 216.590 -26.610 217.690 -26.560 ;
        RECT 216.590 -26.650 217.030 -26.610 ;
        RECT 199.010 -27.220 199.460 -27.140 ;
        RECT 197.160 -27.460 199.460 -27.220 ;
        RECT 197.160 -27.560 197.610 -27.460 ;
        RECT 199.010 -27.560 199.460 -27.460 ;
        RECT 200.410 -27.220 200.860 -27.110 ;
        RECT 202.260 -27.220 202.710 -27.110 ;
        RECT 200.410 -27.460 202.710 -27.220 ;
        RECT 200.410 -27.530 200.860 -27.460 ;
        RECT 183.660 -28.090 184.110 -28.040 ;
        RECT 182.020 -28.380 184.110 -28.090 ;
        RECT 182.020 -28.430 182.470 -28.380 ;
        RECT 165.270 -29.010 165.720 -28.940 ;
        RECT 163.420 -29.250 165.720 -29.010 ;
        RECT 163.420 -29.360 163.870 -29.250 ;
        RECT 165.270 -29.360 165.720 -29.250 ;
        RECT 166.670 -29.010 167.120 -28.910 ;
        RECT 168.520 -29.010 168.970 -28.910 ;
        RECT 166.670 -29.250 168.970 -29.010 ;
        RECT 166.670 -29.330 167.120 -29.250 ;
        RECT 147.180 -29.910 148.710 -29.700 ;
        RECT 149.090 -29.910 149.540 -29.820 ;
        RECT 149.920 -29.910 151.450 -29.700 ;
        RECT 160.680 -29.700 161.130 -29.420 ;
        RECT 164.500 -29.700 164.950 -29.420 ;
        RECT 167.720 -29.690 168.130 -29.250 ;
        RECT 168.520 -29.360 168.970 -29.250 ;
        RECT 170.160 -29.010 170.610 -28.910 ;
        RECT 172.010 -29.010 172.460 -28.910 ;
        RECT 170.160 -29.250 172.460 -29.010 ;
        RECT 170.160 -29.360 170.610 -29.250 ;
        RECT 171.000 -29.690 171.410 -29.250 ;
        RECT 172.010 -29.330 172.460 -29.250 ;
        RECT 173.410 -29.010 173.860 -28.940 ;
        RECT 174.460 -29.010 174.870 -28.580 ;
        RECT 175.260 -29.010 175.710 -28.910 ;
        RECT 173.410 -29.250 175.710 -29.010 ;
        RECT 173.410 -29.360 173.860 -29.250 ;
        RECT 175.260 -29.360 175.710 -29.250 ;
        RECT 176.920 -29.010 177.370 -28.910 ;
        RECT 177.760 -29.010 178.170 -28.580 ;
        RECT 180.920 -28.650 182.470 -28.430 ;
        RECT 182.850 -28.440 183.280 -28.380 ;
        RECT 183.660 -28.430 184.110 -28.380 ;
        RECT 184.710 -28.430 185.210 -28.040 ;
        RECT 183.660 -28.650 185.210 -28.430 ;
        RECT 194.420 -28.040 195.970 -27.820 ;
        RECT 194.420 -28.430 194.920 -28.040 ;
        RECT 195.520 -28.090 195.970 -28.040 ;
        RECT 196.350 -28.090 196.780 -28.030 ;
        RECT 197.160 -28.040 198.710 -27.820 ;
        RECT 201.460 -27.890 201.870 -27.460 ;
        RECT 202.260 -27.560 202.710 -27.460 ;
        RECT 203.920 -27.220 204.370 -27.110 ;
        RECT 205.770 -27.220 206.220 -27.110 ;
        RECT 203.920 -27.460 206.220 -27.220 ;
        RECT 203.920 -27.560 204.370 -27.460 ;
        RECT 204.760 -27.890 205.170 -27.460 ;
        RECT 205.770 -27.530 206.220 -27.460 ;
        RECT 207.170 -27.220 207.620 -27.140 ;
        RECT 208.220 -27.220 208.630 -26.780 ;
        RECT 209.020 -27.220 209.470 -27.110 ;
        RECT 207.170 -27.460 209.470 -27.220 ;
        RECT 207.170 -27.560 207.620 -27.460 ;
        RECT 209.020 -27.560 209.470 -27.460 ;
        RECT 210.660 -27.220 211.110 -27.110 ;
        RECT 211.500 -27.220 211.910 -26.780 ;
        RECT 214.680 -27.050 215.130 -26.770 ;
        RECT 212.510 -27.220 212.960 -27.140 ;
        RECT 210.660 -27.460 212.960 -27.220 ;
        RECT 210.660 -27.560 211.110 -27.460 ;
        RECT 212.510 -27.560 212.960 -27.460 ;
        RECT 213.910 -27.220 214.360 -27.110 ;
        RECT 215.760 -27.220 216.210 -27.110 ;
        RECT 213.910 -27.460 216.210 -27.220 ;
        RECT 213.910 -27.530 214.360 -27.460 ;
        RECT 197.160 -28.090 197.610 -28.040 ;
        RECT 195.520 -28.380 197.610 -28.090 ;
        RECT 195.520 -28.430 195.970 -28.380 ;
        RECT 178.770 -29.010 179.220 -28.940 ;
        RECT 176.920 -29.250 179.220 -29.010 ;
        RECT 176.920 -29.360 177.370 -29.250 ;
        RECT 178.770 -29.360 179.220 -29.250 ;
        RECT 180.170 -29.010 180.620 -28.910 ;
        RECT 182.020 -29.010 182.470 -28.910 ;
        RECT 180.170 -29.250 182.470 -29.010 ;
        RECT 180.170 -29.330 180.620 -29.250 ;
        RECT 160.680 -29.910 162.210 -29.700 ;
        RECT 162.590 -29.910 163.040 -29.820 ;
        RECT 163.420 -29.910 164.950 -29.700 ;
        RECT 174.180 -29.700 174.630 -29.420 ;
        RECT 178.000 -29.700 178.450 -29.420 ;
        RECT 181.220 -29.690 181.630 -29.250 ;
        RECT 182.020 -29.360 182.470 -29.250 ;
        RECT 183.660 -29.010 184.110 -28.910 ;
        RECT 185.510 -29.010 185.960 -28.910 ;
        RECT 183.660 -29.250 185.960 -29.010 ;
        RECT 183.660 -29.360 184.110 -29.250 ;
        RECT 184.500 -29.690 184.910 -29.250 ;
        RECT 185.510 -29.330 185.960 -29.250 ;
        RECT 186.910 -29.010 187.360 -28.940 ;
        RECT 187.960 -29.010 188.370 -28.580 ;
        RECT 188.760 -29.010 189.210 -28.910 ;
        RECT 186.910 -29.250 189.210 -29.010 ;
        RECT 186.910 -29.360 187.360 -29.250 ;
        RECT 188.760 -29.360 189.210 -29.250 ;
        RECT 190.420 -29.010 190.870 -28.910 ;
        RECT 191.260 -29.010 191.670 -28.580 ;
        RECT 194.420 -28.650 195.970 -28.430 ;
        RECT 196.350 -28.440 196.780 -28.380 ;
        RECT 197.160 -28.430 197.610 -28.380 ;
        RECT 198.210 -28.430 198.710 -28.040 ;
        RECT 197.160 -28.650 198.710 -28.430 ;
        RECT 207.920 -28.040 209.470 -27.820 ;
        RECT 207.920 -28.430 208.420 -28.040 ;
        RECT 209.020 -28.090 209.470 -28.040 ;
        RECT 209.850 -28.090 210.280 -28.030 ;
        RECT 210.660 -28.040 212.210 -27.820 ;
        RECT 214.960 -27.890 215.370 -27.460 ;
        RECT 215.760 -27.560 216.210 -27.460 ;
        RECT 210.660 -28.090 211.110 -28.040 ;
        RECT 209.020 -28.380 211.110 -28.090 ;
        RECT 209.020 -28.430 209.470 -28.380 ;
        RECT 192.270 -29.010 192.720 -28.940 ;
        RECT 190.420 -29.250 192.720 -29.010 ;
        RECT 190.420 -29.360 190.870 -29.250 ;
        RECT 192.270 -29.360 192.720 -29.250 ;
        RECT 193.670 -29.010 194.120 -28.910 ;
        RECT 195.520 -29.010 195.970 -28.910 ;
        RECT 193.670 -29.250 195.970 -29.010 ;
        RECT 193.670 -29.330 194.120 -29.250 ;
        RECT 174.180 -29.910 175.710 -29.700 ;
        RECT 176.090 -29.910 176.540 -29.820 ;
        RECT 176.920 -29.910 178.450 -29.700 ;
        RECT 187.680 -29.700 188.130 -29.420 ;
        RECT 191.500 -29.700 191.950 -29.420 ;
        RECT 194.720 -29.690 195.130 -29.250 ;
        RECT 195.520 -29.360 195.970 -29.250 ;
        RECT 197.160 -29.010 197.610 -28.910 ;
        RECT 199.010 -29.010 199.460 -28.910 ;
        RECT 197.160 -29.250 199.460 -29.010 ;
        RECT 197.160 -29.360 197.610 -29.250 ;
        RECT 198.000 -29.690 198.410 -29.250 ;
        RECT 199.010 -29.330 199.460 -29.250 ;
        RECT 200.410 -29.010 200.860 -28.940 ;
        RECT 201.460 -29.010 201.870 -28.580 ;
        RECT 202.260 -29.010 202.710 -28.910 ;
        RECT 200.410 -29.250 202.710 -29.010 ;
        RECT 200.410 -29.360 200.860 -29.250 ;
        RECT 202.260 -29.360 202.710 -29.250 ;
        RECT 203.920 -29.010 204.370 -28.910 ;
        RECT 204.760 -29.010 205.170 -28.580 ;
        RECT 207.920 -28.650 209.470 -28.430 ;
        RECT 209.850 -28.440 210.280 -28.380 ;
        RECT 210.660 -28.430 211.110 -28.380 ;
        RECT 211.710 -28.430 212.210 -28.040 ;
        RECT 210.660 -28.650 212.210 -28.430 ;
        RECT 205.770 -29.010 206.220 -28.940 ;
        RECT 203.920 -29.250 206.220 -29.010 ;
        RECT 203.920 -29.360 204.370 -29.250 ;
        RECT 205.770 -29.360 206.220 -29.250 ;
        RECT 207.170 -29.010 207.620 -28.910 ;
        RECT 209.020 -29.010 209.470 -28.910 ;
        RECT 207.170 -29.250 209.470 -29.010 ;
        RECT 207.170 -29.330 207.620 -29.250 ;
        RECT 187.680 -29.910 189.210 -29.700 ;
        RECT 189.590 -29.910 190.040 -29.820 ;
        RECT 190.420 -29.910 191.950 -29.700 ;
        RECT 201.180 -29.700 201.630 -29.420 ;
        RECT 205.000 -29.700 205.450 -29.420 ;
        RECT 208.220 -29.690 208.630 -29.250 ;
        RECT 209.020 -29.360 209.470 -29.250 ;
        RECT 210.660 -29.010 211.110 -28.910 ;
        RECT 212.510 -29.010 212.960 -28.910 ;
        RECT 210.660 -29.250 212.960 -29.010 ;
        RECT 210.660 -29.360 211.110 -29.250 ;
        RECT 211.500 -29.690 211.910 -29.250 ;
        RECT 212.510 -29.330 212.960 -29.250 ;
        RECT 213.910 -29.010 214.360 -28.940 ;
        RECT 214.960 -29.010 215.370 -28.580 ;
        RECT 215.760 -29.010 216.210 -28.910 ;
        RECT 213.910 -29.250 216.210 -29.010 ;
        RECT 213.910 -29.360 214.360 -29.250 ;
        RECT 215.760 -29.360 216.210 -29.250 ;
        RECT 201.180 -29.910 202.710 -29.700 ;
        RECT 203.090 -29.910 203.540 -29.820 ;
        RECT 203.920 -29.910 205.450 -29.700 ;
        RECT 214.680 -29.700 215.130 -29.420 ;
        RECT 214.680 -29.910 216.210 -29.700 ;
        RECT 216.590 -29.910 217.030 -29.820 ;
        RECT 13.260 -30.170 15.370 -29.910 ;
        RECT 26.760 -30.170 28.870 -29.910 ;
        RECT 40.260 -30.170 42.370 -29.910 ;
        RECT 53.760 -30.170 55.870 -29.910 ;
        RECT 67.260 -30.170 69.370 -29.910 ;
        RECT 80.760 -30.170 82.870 -29.910 ;
        RECT 94.260 -30.170 96.370 -29.910 ;
        RECT 107.760 -30.170 109.870 -29.910 ;
        RECT 121.260 -30.170 123.370 -29.910 ;
        RECT 134.760 -30.170 136.870 -29.910 ;
        RECT 148.260 -30.170 150.370 -29.910 ;
        RECT 161.760 -30.170 163.870 -29.910 ;
        RECT 175.260 -30.170 177.370 -29.910 ;
        RECT 188.760 -30.170 190.870 -29.910 ;
        RECT 202.260 -30.170 204.370 -29.910 ;
        RECT 215.760 -29.920 217.030 -29.910 ;
        RECT 215.760 -30.110 217.240 -29.920 ;
        RECT 215.760 -30.170 217.030 -30.110 ;
        RECT 12.180 -30.380 13.710 -30.170 ;
        RECT 14.090 -30.260 14.540 -30.170 ;
        RECT 14.920 -30.380 16.450 -30.170 ;
        RECT 1.420 -30.830 1.870 -30.720 ;
        RECT 3.270 -30.830 3.720 -30.720 ;
        RECT 1.420 -31.070 3.720 -30.830 ;
        RECT 1.420 -31.170 1.870 -31.070 ;
        RECT 2.260 -31.500 2.670 -31.070 ;
        RECT 3.270 -31.140 3.720 -31.070 ;
        RECT 4.670 -30.830 5.120 -30.750 ;
        RECT 5.720 -30.830 6.130 -30.390 ;
        RECT 6.520 -30.830 6.970 -30.720 ;
        RECT 4.670 -31.070 6.970 -30.830 ;
        RECT 4.670 -31.170 5.120 -31.070 ;
        RECT 6.520 -31.170 6.970 -31.070 ;
        RECT 8.160 -30.830 8.610 -30.720 ;
        RECT 9.000 -30.830 9.410 -30.390 ;
        RECT 12.180 -30.660 12.630 -30.380 ;
        RECT 16.000 -30.660 16.450 -30.380 ;
        RECT 25.680 -30.380 27.210 -30.170 ;
        RECT 27.590 -30.260 28.040 -30.170 ;
        RECT 28.420 -30.380 29.950 -30.170 ;
        RECT 10.010 -30.830 10.460 -30.750 ;
        RECT 8.160 -31.070 10.460 -30.830 ;
        RECT 8.160 -31.170 8.610 -31.070 ;
        RECT 10.010 -31.170 10.460 -31.070 ;
        RECT 11.410 -30.830 11.860 -30.720 ;
        RECT 13.260 -30.830 13.710 -30.720 ;
        RECT 11.410 -31.070 13.710 -30.830 ;
        RECT 11.410 -31.140 11.860 -31.070 ;
        RECT 5.420 -31.650 6.970 -31.430 ;
        RECT 5.420 -32.040 5.920 -31.650 ;
        RECT 6.520 -31.700 6.970 -31.650 ;
        RECT 7.350 -31.700 7.780 -31.640 ;
        RECT 8.160 -31.650 9.710 -31.430 ;
        RECT 12.460 -31.500 12.870 -31.070 ;
        RECT 13.260 -31.170 13.710 -31.070 ;
        RECT 14.920 -30.830 15.370 -30.720 ;
        RECT 16.770 -30.830 17.220 -30.720 ;
        RECT 14.920 -31.070 17.220 -30.830 ;
        RECT 14.920 -31.170 15.370 -31.070 ;
        RECT 15.760 -31.500 16.170 -31.070 ;
        RECT 16.770 -31.140 17.220 -31.070 ;
        RECT 18.170 -30.830 18.620 -30.750 ;
        RECT 19.220 -30.830 19.630 -30.390 ;
        RECT 20.020 -30.830 20.470 -30.720 ;
        RECT 18.170 -31.070 20.470 -30.830 ;
        RECT 18.170 -31.170 18.620 -31.070 ;
        RECT 20.020 -31.170 20.470 -31.070 ;
        RECT 21.660 -30.830 22.110 -30.720 ;
        RECT 22.500 -30.830 22.910 -30.390 ;
        RECT 25.680 -30.660 26.130 -30.380 ;
        RECT 29.500 -30.660 29.950 -30.380 ;
        RECT 39.180 -30.380 40.710 -30.170 ;
        RECT 41.090 -30.260 41.540 -30.170 ;
        RECT 41.920 -30.380 43.450 -30.170 ;
        RECT 23.510 -30.830 23.960 -30.750 ;
        RECT 21.660 -31.070 23.960 -30.830 ;
        RECT 21.660 -31.170 22.110 -31.070 ;
        RECT 23.510 -31.170 23.960 -31.070 ;
        RECT 24.910 -30.830 25.360 -30.720 ;
        RECT 26.760 -30.830 27.210 -30.720 ;
        RECT 24.910 -31.070 27.210 -30.830 ;
        RECT 24.910 -31.140 25.360 -31.070 ;
        RECT 8.160 -31.700 8.610 -31.650 ;
        RECT 6.520 -31.990 8.610 -31.700 ;
        RECT 6.520 -32.040 6.970 -31.990 ;
        RECT 1.420 -32.620 1.870 -32.520 ;
        RECT 2.260 -32.620 2.670 -32.190 ;
        RECT 5.420 -32.260 6.970 -32.040 ;
        RECT 7.350 -32.050 7.780 -31.990 ;
        RECT 8.160 -32.040 8.610 -31.990 ;
        RECT 9.210 -32.040 9.710 -31.650 ;
        RECT 8.160 -32.260 9.710 -32.040 ;
        RECT 18.920 -31.650 20.470 -31.430 ;
        RECT 18.920 -32.040 19.420 -31.650 ;
        RECT 20.020 -31.700 20.470 -31.650 ;
        RECT 20.850 -31.700 21.280 -31.640 ;
        RECT 21.660 -31.650 23.210 -31.430 ;
        RECT 25.960 -31.500 26.370 -31.070 ;
        RECT 26.760 -31.170 27.210 -31.070 ;
        RECT 28.420 -30.830 28.870 -30.720 ;
        RECT 30.270 -30.830 30.720 -30.720 ;
        RECT 28.420 -31.070 30.720 -30.830 ;
        RECT 28.420 -31.170 28.870 -31.070 ;
        RECT 29.260 -31.500 29.670 -31.070 ;
        RECT 30.270 -31.140 30.720 -31.070 ;
        RECT 31.670 -30.830 32.120 -30.750 ;
        RECT 32.720 -30.830 33.130 -30.390 ;
        RECT 33.520 -30.830 33.970 -30.720 ;
        RECT 31.670 -31.070 33.970 -30.830 ;
        RECT 31.670 -31.170 32.120 -31.070 ;
        RECT 33.520 -31.170 33.970 -31.070 ;
        RECT 35.160 -30.830 35.610 -30.720 ;
        RECT 36.000 -30.830 36.410 -30.390 ;
        RECT 39.180 -30.660 39.630 -30.380 ;
        RECT 43.000 -30.660 43.450 -30.380 ;
        RECT 52.680 -30.380 54.210 -30.170 ;
        RECT 54.590 -30.260 55.040 -30.170 ;
        RECT 55.420 -30.380 56.950 -30.170 ;
        RECT 37.010 -30.830 37.460 -30.750 ;
        RECT 35.160 -31.070 37.460 -30.830 ;
        RECT 35.160 -31.170 35.610 -31.070 ;
        RECT 37.010 -31.170 37.460 -31.070 ;
        RECT 38.410 -30.830 38.860 -30.720 ;
        RECT 40.260 -30.830 40.710 -30.720 ;
        RECT 38.410 -31.070 40.710 -30.830 ;
        RECT 38.410 -31.140 38.860 -31.070 ;
        RECT 21.660 -31.700 22.110 -31.650 ;
        RECT 20.020 -31.990 22.110 -31.700 ;
        RECT 20.020 -32.040 20.470 -31.990 ;
        RECT 3.270 -32.620 3.720 -32.550 ;
        RECT 1.420 -32.860 3.720 -32.620 ;
        RECT 1.420 -32.970 1.870 -32.860 ;
        RECT 3.270 -32.970 3.720 -32.860 ;
        RECT 4.670 -32.620 5.120 -32.520 ;
        RECT 6.520 -32.620 6.970 -32.520 ;
        RECT 4.670 -32.860 6.970 -32.620 ;
        RECT 4.670 -32.940 5.120 -32.860 ;
        RECT 5.720 -33.300 6.130 -32.860 ;
        RECT 6.520 -32.970 6.970 -32.860 ;
        RECT 8.160 -32.620 8.610 -32.520 ;
        RECT 10.010 -32.620 10.460 -32.520 ;
        RECT 8.160 -32.860 10.460 -32.620 ;
        RECT 8.160 -32.970 8.610 -32.860 ;
        RECT 9.000 -33.300 9.410 -32.860 ;
        RECT 10.010 -32.940 10.460 -32.860 ;
        RECT 11.410 -32.620 11.860 -32.550 ;
        RECT 12.460 -32.620 12.870 -32.190 ;
        RECT 13.260 -32.620 13.710 -32.520 ;
        RECT 11.410 -32.860 13.710 -32.620 ;
        RECT 11.410 -32.970 11.860 -32.860 ;
        RECT 13.260 -32.970 13.710 -32.860 ;
        RECT 14.920 -32.620 15.370 -32.520 ;
        RECT 15.760 -32.620 16.170 -32.190 ;
        RECT 18.920 -32.260 20.470 -32.040 ;
        RECT 20.850 -32.050 21.280 -31.990 ;
        RECT 21.660 -32.040 22.110 -31.990 ;
        RECT 22.710 -32.040 23.210 -31.650 ;
        RECT 21.660 -32.260 23.210 -32.040 ;
        RECT 32.420 -31.650 33.970 -31.430 ;
        RECT 32.420 -32.040 32.920 -31.650 ;
        RECT 33.520 -31.700 33.970 -31.650 ;
        RECT 34.350 -31.700 34.780 -31.640 ;
        RECT 35.160 -31.650 36.710 -31.430 ;
        RECT 39.460 -31.500 39.870 -31.070 ;
        RECT 40.260 -31.170 40.710 -31.070 ;
        RECT 41.920 -30.830 42.370 -30.720 ;
        RECT 43.770 -30.830 44.220 -30.720 ;
        RECT 41.920 -31.070 44.220 -30.830 ;
        RECT 41.920 -31.170 42.370 -31.070 ;
        RECT 42.760 -31.500 43.170 -31.070 ;
        RECT 43.770 -31.140 44.220 -31.070 ;
        RECT 45.170 -30.830 45.620 -30.750 ;
        RECT 46.220 -30.830 46.630 -30.390 ;
        RECT 47.020 -30.830 47.470 -30.720 ;
        RECT 45.170 -31.070 47.470 -30.830 ;
        RECT 45.170 -31.170 45.620 -31.070 ;
        RECT 47.020 -31.170 47.470 -31.070 ;
        RECT 48.660 -30.830 49.110 -30.720 ;
        RECT 49.500 -30.830 49.910 -30.390 ;
        RECT 52.680 -30.660 53.130 -30.380 ;
        RECT 56.500 -30.660 56.950 -30.380 ;
        RECT 66.180 -30.380 67.710 -30.170 ;
        RECT 68.090 -30.260 68.540 -30.170 ;
        RECT 68.920 -30.380 70.450 -30.170 ;
        RECT 50.510 -30.830 50.960 -30.750 ;
        RECT 48.660 -31.070 50.960 -30.830 ;
        RECT 48.660 -31.170 49.110 -31.070 ;
        RECT 50.510 -31.170 50.960 -31.070 ;
        RECT 51.910 -30.830 52.360 -30.720 ;
        RECT 53.760 -30.830 54.210 -30.720 ;
        RECT 51.910 -31.070 54.210 -30.830 ;
        RECT 51.910 -31.140 52.360 -31.070 ;
        RECT 35.160 -31.700 35.610 -31.650 ;
        RECT 33.520 -31.990 35.610 -31.700 ;
        RECT 33.520 -32.040 33.970 -31.990 ;
        RECT 16.770 -32.620 17.220 -32.550 ;
        RECT 14.920 -32.860 17.220 -32.620 ;
        RECT 14.920 -32.970 15.370 -32.860 ;
        RECT 16.770 -32.970 17.220 -32.860 ;
        RECT 18.170 -32.620 18.620 -32.520 ;
        RECT 20.020 -32.620 20.470 -32.520 ;
        RECT 18.170 -32.860 20.470 -32.620 ;
        RECT 18.170 -32.940 18.620 -32.860 ;
        RECT 12.180 -33.310 12.630 -33.030 ;
        RECT 16.000 -33.310 16.450 -33.030 ;
        RECT 19.220 -33.300 19.630 -32.860 ;
        RECT 20.020 -32.970 20.470 -32.860 ;
        RECT 21.660 -32.620 22.110 -32.520 ;
        RECT 23.510 -32.620 23.960 -32.520 ;
        RECT 21.660 -32.860 23.960 -32.620 ;
        RECT 21.660 -32.970 22.110 -32.860 ;
        RECT 22.500 -33.300 22.910 -32.860 ;
        RECT 23.510 -32.940 23.960 -32.860 ;
        RECT 24.910 -32.620 25.360 -32.550 ;
        RECT 25.960 -32.620 26.370 -32.190 ;
        RECT 26.760 -32.620 27.210 -32.520 ;
        RECT 24.910 -32.860 27.210 -32.620 ;
        RECT 24.910 -32.970 25.360 -32.860 ;
        RECT 26.760 -32.970 27.210 -32.860 ;
        RECT 28.420 -32.620 28.870 -32.520 ;
        RECT 29.260 -32.620 29.670 -32.190 ;
        RECT 32.420 -32.260 33.970 -32.040 ;
        RECT 34.350 -32.050 34.780 -31.990 ;
        RECT 35.160 -32.040 35.610 -31.990 ;
        RECT 36.210 -32.040 36.710 -31.650 ;
        RECT 35.160 -32.260 36.710 -32.040 ;
        RECT 45.920 -31.650 47.470 -31.430 ;
        RECT 45.920 -32.040 46.420 -31.650 ;
        RECT 47.020 -31.700 47.470 -31.650 ;
        RECT 47.850 -31.700 48.280 -31.640 ;
        RECT 48.660 -31.650 50.210 -31.430 ;
        RECT 52.960 -31.500 53.370 -31.070 ;
        RECT 53.760 -31.170 54.210 -31.070 ;
        RECT 55.420 -30.830 55.870 -30.720 ;
        RECT 57.270 -30.830 57.720 -30.720 ;
        RECT 55.420 -31.070 57.720 -30.830 ;
        RECT 55.420 -31.170 55.870 -31.070 ;
        RECT 56.260 -31.500 56.670 -31.070 ;
        RECT 57.270 -31.140 57.720 -31.070 ;
        RECT 58.670 -30.830 59.120 -30.750 ;
        RECT 59.720 -30.830 60.130 -30.390 ;
        RECT 60.520 -30.830 60.970 -30.720 ;
        RECT 58.670 -31.070 60.970 -30.830 ;
        RECT 58.670 -31.170 59.120 -31.070 ;
        RECT 60.520 -31.170 60.970 -31.070 ;
        RECT 62.160 -30.830 62.610 -30.720 ;
        RECT 63.000 -30.830 63.410 -30.390 ;
        RECT 66.180 -30.660 66.630 -30.380 ;
        RECT 70.000 -30.660 70.450 -30.380 ;
        RECT 79.680 -30.380 81.210 -30.170 ;
        RECT 81.590 -30.260 82.040 -30.170 ;
        RECT 82.420 -30.380 83.950 -30.170 ;
        RECT 64.010 -30.830 64.460 -30.750 ;
        RECT 62.160 -31.070 64.460 -30.830 ;
        RECT 62.160 -31.170 62.610 -31.070 ;
        RECT 64.010 -31.170 64.460 -31.070 ;
        RECT 65.410 -30.830 65.860 -30.720 ;
        RECT 67.260 -30.830 67.710 -30.720 ;
        RECT 65.410 -31.070 67.710 -30.830 ;
        RECT 65.410 -31.140 65.860 -31.070 ;
        RECT 48.660 -31.700 49.110 -31.650 ;
        RECT 47.020 -31.990 49.110 -31.700 ;
        RECT 47.020 -32.040 47.470 -31.990 ;
        RECT 30.270 -32.620 30.720 -32.550 ;
        RECT 28.420 -32.860 30.720 -32.620 ;
        RECT 28.420 -32.970 28.870 -32.860 ;
        RECT 30.270 -32.970 30.720 -32.860 ;
        RECT 31.670 -32.620 32.120 -32.520 ;
        RECT 33.520 -32.620 33.970 -32.520 ;
        RECT 31.670 -32.860 33.970 -32.620 ;
        RECT 31.670 -32.940 32.120 -32.860 ;
        RECT 12.180 -33.520 13.710 -33.310 ;
        RECT 14.090 -33.520 14.540 -33.430 ;
        RECT 14.920 -33.520 16.450 -33.310 ;
        RECT 25.680 -33.310 26.130 -33.030 ;
        RECT 29.500 -33.310 29.950 -33.030 ;
        RECT 32.720 -33.300 33.130 -32.860 ;
        RECT 33.520 -32.970 33.970 -32.860 ;
        RECT 35.160 -32.620 35.610 -32.520 ;
        RECT 37.010 -32.620 37.460 -32.520 ;
        RECT 35.160 -32.860 37.460 -32.620 ;
        RECT 35.160 -32.970 35.610 -32.860 ;
        RECT 36.000 -33.300 36.410 -32.860 ;
        RECT 37.010 -32.940 37.460 -32.860 ;
        RECT 38.410 -32.620 38.860 -32.550 ;
        RECT 39.460 -32.620 39.870 -32.190 ;
        RECT 40.260 -32.620 40.710 -32.520 ;
        RECT 38.410 -32.860 40.710 -32.620 ;
        RECT 38.410 -32.970 38.860 -32.860 ;
        RECT 40.260 -32.970 40.710 -32.860 ;
        RECT 41.920 -32.620 42.370 -32.520 ;
        RECT 42.760 -32.620 43.170 -32.190 ;
        RECT 45.920 -32.260 47.470 -32.040 ;
        RECT 47.850 -32.050 48.280 -31.990 ;
        RECT 48.660 -32.040 49.110 -31.990 ;
        RECT 49.710 -32.040 50.210 -31.650 ;
        RECT 48.660 -32.260 50.210 -32.040 ;
        RECT 59.420 -31.650 60.970 -31.430 ;
        RECT 59.420 -32.040 59.920 -31.650 ;
        RECT 60.520 -31.700 60.970 -31.650 ;
        RECT 61.350 -31.700 61.780 -31.640 ;
        RECT 62.160 -31.650 63.710 -31.430 ;
        RECT 66.460 -31.500 66.870 -31.070 ;
        RECT 67.260 -31.170 67.710 -31.070 ;
        RECT 68.920 -30.830 69.370 -30.720 ;
        RECT 70.770 -30.830 71.220 -30.720 ;
        RECT 68.920 -31.070 71.220 -30.830 ;
        RECT 68.920 -31.170 69.370 -31.070 ;
        RECT 69.760 -31.500 70.170 -31.070 ;
        RECT 70.770 -31.140 71.220 -31.070 ;
        RECT 72.170 -30.830 72.620 -30.750 ;
        RECT 73.220 -30.830 73.630 -30.390 ;
        RECT 74.020 -30.830 74.470 -30.720 ;
        RECT 72.170 -31.070 74.470 -30.830 ;
        RECT 72.170 -31.170 72.620 -31.070 ;
        RECT 74.020 -31.170 74.470 -31.070 ;
        RECT 75.660 -30.830 76.110 -30.720 ;
        RECT 76.500 -30.830 76.910 -30.390 ;
        RECT 79.680 -30.660 80.130 -30.380 ;
        RECT 83.500 -30.660 83.950 -30.380 ;
        RECT 93.180 -30.380 94.710 -30.170 ;
        RECT 95.090 -30.260 95.540 -30.170 ;
        RECT 95.920 -30.380 97.450 -30.170 ;
        RECT 77.510 -30.830 77.960 -30.750 ;
        RECT 75.660 -31.070 77.960 -30.830 ;
        RECT 75.660 -31.170 76.110 -31.070 ;
        RECT 77.510 -31.170 77.960 -31.070 ;
        RECT 78.910 -30.830 79.360 -30.720 ;
        RECT 80.760 -30.830 81.210 -30.720 ;
        RECT 78.910 -31.070 81.210 -30.830 ;
        RECT 78.910 -31.140 79.360 -31.070 ;
        RECT 62.160 -31.700 62.610 -31.650 ;
        RECT 60.520 -31.990 62.610 -31.700 ;
        RECT 60.520 -32.040 60.970 -31.990 ;
        RECT 43.770 -32.620 44.220 -32.550 ;
        RECT 41.920 -32.860 44.220 -32.620 ;
        RECT 41.920 -32.970 42.370 -32.860 ;
        RECT 43.770 -32.970 44.220 -32.860 ;
        RECT 45.170 -32.620 45.620 -32.520 ;
        RECT 47.020 -32.620 47.470 -32.520 ;
        RECT 45.170 -32.860 47.470 -32.620 ;
        RECT 45.170 -32.940 45.620 -32.860 ;
        RECT 25.680 -33.520 27.210 -33.310 ;
        RECT 27.590 -33.520 28.040 -33.430 ;
        RECT 28.420 -33.520 29.950 -33.310 ;
        RECT 39.180 -33.310 39.630 -33.030 ;
        RECT 43.000 -33.310 43.450 -33.030 ;
        RECT 46.220 -33.300 46.630 -32.860 ;
        RECT 47.020 -32.970 47.470 -32.860 ;
        RECT 48.660 -32.620 49.110 -32.520 ;
        RECT 50.510 -32.620 50.960 -32.520 ;
        RECT 48.660 -32.860 50.960 -32.620 ;
        RECT 48.660 -32.970 49.110 -32.860 ;
        RECT 49.500 -33.300 49.910 -32.860 ;
        RECT 50.510 -32.940 50.960 -32.860 ;
        RECT 51.910 -32.620 52.360 -32.550 ;
        RECT 52.960 -32.620 53.370 -32.190 ;
        RECT 53.760 -32.620 54.210 -32.520 ;
        RECT 51.910 -32.860 54.210 -32.620 ;
        RECT 51.910 -32.970 52.360 -32.860 ;
        RECT 53.760 -32.970 54.210 -32.860 ;
        RECT 55.420 -32.620 55.870 -32.520 ;
        RECT 56.260 -32.620 56.670 -32.190 ;
        RECT 59.420 -32.260 60.970 -32.040 ;
        RECT 61.350 -32.050 61.780 -31.990 ;
        RECT 62.160 -32.040 62.610 -31.990 ;
        RECT 63.210 -32.040 63.710 -31.650 ;
        RECT 62.160 -32.260 63.710 -32.040 ;
        RECT 72.920 -31.650 74.470 -31.430 ;
        RECT 72.920 -32.040 73.420 -31.650 ;
        RECT 74.020 -31.700 74.470 -31.650 ;
        RECT 74.850 -31.700 75.280 -31.640 ;
        RECT 75.660 -31.650 77.210 -31.430 ;
        RECT 79.960 -31.500 80.370 -31.070 ;
        RECT 80.760 -31.170 81.210 -31.070 ;
        RECT 82.420 -30.830 82.870 -30.720 ;
        RECT 84.270 -30.830 84.720 -30.720 ;
        RECT 82.420 -31.070 84.720 -30.830 ;
        RECT 82.420 -31.170 82.870 -31.070 ;
        RECT 83.260 -31.500 83.670 -31.070 ;
        RECT 84.270 -31.140 84.720 -31.070 ;
        RECT 85.670 -30.830 86.120 -30.750 ;
        RECT 86.720 -30.830 87.130 -30.390 ;
        RECT 87.520 -30.830 87.970 -30.720 ;
        RECT 85.670 -31.070 87.970 -30.830 ;
        RECT 85.670 -31.170 86.120 -31.070 ;
        RECT 87.520 -31.170 87.970 -31.070 ;
        RECT 89.160 -30.830 89.610 -30.720 ;
        RECT 90.000 -30.830 90.410 -30.390 ;
        RECT 93.180 -30.660 93.630 -30.380 ;
        RECT 97.000 -30.660 97.450 -30.380 ;
        RECT 106.680 -30.380 108.210 -30.170 ;
        RECT 108.590 -30.260 109.040 -30.170 ;
        RECT 109.420 -30.380 110.950 -30.170 ;
        RECT 91.010 -30.830 91.460 -30.750 ;
        RECT 89.160 -31.070 91.460 -30.830 ;
        RECT 89.160 -31.170 89.610 -31.070 ;
        RECT 91.010 -31.170 91.460 -31.070 ;
        RECT 92.410 -30.830 92.860 -30.720 ;
        RECT 94.260 -30.830 94.710 -30.720 ;
        RECT 92.410 -31.070 94.710 -30.830 ;
        RECT 92.410 -31.140 92.860 -31.070 ;
        RECT 75.660 -31.700 76.110 -31.650 ;
        RECT 74.020 -31.990 76.110 -31.700 ;
        RECT 74.020 -32.040 74.470 -31.990 ;
        RECT 57.270 -32.620 57.720 -32.550 ;
        RECT 55.420 -32.860 57.720 -32.620 ;
        RECT 55.420 -32.970 55.870 -32.860 ;
        RECT 57.270 -32.970 57.720 -32.860 ;
        RECT 58.670 -32.620 59.120 -32.520 ;
        RECT 60.520 -32.620 60.970 -32.520 ;
        RECT 58.670 -32.860 60.970 -32.620 ;
        RECT 58.670 -32.940 59.120 -32.860 ;
        RECT 39.180 -33.520 40.710 -33.310 ;
        RECT 41.090 -33.520 41.540 -33.430 ;
        RECT 41.920 -33.520 43.450 -33.310 ;
        RECT 52.680 -33.310 53.130 -33.030 ;
        RECT 56.500 -33.310 56.950 -33.030 ;
        RECT 59.720 -33.300 60.130 -32.860 ;
        RECT 60.520 -32.970 60.970 -32.860 ;
        RECT 62.160 -32.620 62.610 -32.520 ;
        RECT 64.010 -32.620 64.460 -32.520 ;
        RECT 62.160 -32.860 64.460 -32.620 ;
        RECT 62.160 -32.970 62.610 -32.860 ;
        RECT 63.000 -33.300 63.410 -32.860 ;
        RECT 64.010 -32.940 64.460 -32.860 ;
        RECT 65.410 -32.620 65.860 -32.550 ;
        RECT 66.460 -32.620 66.870 -32.190 ;
        RECT 67.260 -32.620 67.710 -32.520 ;
        RECT 65.410 -32.860 67.710 -32.620 ;
        RECT 65.410 -32.970 65.860 -32.860 ;
        RECT 67.260 -32.970 67.710 -32.860 ;
        RECT 68.920 -32.620 69.370 -32.520 ;
        RECT 69.760 -32.620 70.170 -32.190 ;
        RECT 72.920 -32.260 74.470 -32.040 ;
        RECT 74.850 -32.050 75.280 -31.990 ;
        RECT 75.660 -32.040 76.110 -31.990 ;
        RECT 76.710 -32.040 77.210 -31.650 ;
        RECT 75.660 -32.260 77.210 -32.040 ;
        RECT 86.420 -31.650 87.970 -31.430 ;
        RECT 86.420 -32.040 86.920 -31.650 ;
        RECT 87.520 -31.700 87.970 -31.650 ;
        RECT 88.350 -31.700 88.780 -31.640 ;
        RECT 89.160 -31.650 90.710 -31.430 ;
        RECT 93.460 -31.500 93.870 -31.070 ;
        RECT 94.260 -31.170 94.710 -31.070 ;
        RECT 95.920 -30.830 96.370 -30.720 ;
        RECT 97.770 -30.830 98.220 -30.720 ;
        RECT 95.920 -31.070 98.220 -30.830 ;
        RECT 95.920 -31.170 96.370 -31.070 ;
        RECT 96.760 -31.500 97.170 -31.070 ;
        RECT 97.770 -31.140 98.220 -31.070 ;
        RECT 99.170 -30.830 99.620 -30.750 ;
        RECT 100.220 -30.830 100.630 -30.390 ;
        RECT 101.020 -30.830 101.470 -30.720 ;
        RECT 99.170 -31.070 101.470 -30.830 ;
        RECT 99.170 -31.170 99.620 -31.070 ;
        RECT 101.020 -31.170 101.470 -31.070 ;
        RECT 102.660 -30.830 103.110 -30.720 ;
        RECT 103.500 -30.830 103.910 -30.390 ;
        RECT 106.680 -30.660 107.130 -30.380 ;
        RECT 110.500 -30.660 110.950 -30.380 ;
        RECT 120.180 -30.380 121.710 -30.170 ;
        RECT 122.090 -30.260 122.540 -30.170 ;
        RECT 122.920 -30.380 124.450 -30.170 ;
        RECT 104.510 -30.830 104.960 -30.750 ;
        RECT 102.660 -31.070 104.960 -30.830 ;
        RECT 102.660 -31.170 103.110 -31.070 ;
        RECT 104.510 -31.170 104.960 -31.070 ;
        RECT 105.910 -30.830 106.360 -30.720 ;
        RECT 107.760 -30.830 108.210 -30.720 ;
        RECT 105.910 -31.070 108.210 -30.830 ;
        RECT 105.910 -31.140 106.360 -31.070 ;
        RECT 89.160 -31.700 89.610 -31.650 ;
        RECT 87.520 -31.990 89.610 -31.700 ;
        RECT 87.520 -32.040 87.970 -31.990 ;
        RECT 70.770 -32.620 71.220 -32.550 ;
        RECT 68.920 -32.860 71.220 -32.620 ;
        RECT 68.920 -32.970 69.370 -32.860 ;
        RECT 70.770 -32.970 71.220 -32.860 ;
        RECT 72.170 -32.620 72.620 -32.520 ;
        RECT 74.020 -32.620 74.470 -32.520 ;
        RECT 72.170 -32.860 74.470 -32.620 ;
        RECT 72.170 -32.940 72.620 -32.860 ;
        RECT 52.680 -33.520 54.210 -33.310 ;
        RECT 54.590 -33.520 55.040 -33.430 ;
        RECT 55.420 -33.520 56.950 -33.310 ;
        RECT 66.180 -33.310 66.630 -33.030 ;
        RECT 70.000 -33.310 70.450 -33.030 ;
        RECT 73.220 -33.300 73.630 -32.860 ;
        RECT 74.020 -32.970 74.470 -32.860 ;
        RECT 75.660 -32.620 76.110 -32.520 ;
        RECT 77.510 -32.620 77.960 -32.520 ;
        RECT 75.660 -32.860 77.960 -32.620 ;
        RECT 75.660 -32.970 76.110 -32.860 ;
        RECT 76.500 -33.300 76.910 -32.860 ;
        RECT 77.510 -32.940 77.960 -32.860 ;
        RECT 78.910 -32.620 79.360 -32.550 ;
        RECT 79.960 -32.620 80.370 -32.190 ;
        RECT 80.760 -32.620 81.210 -32.520 ;
        RECT 78.910 -32.860 81.210 -32.620 ;
        RECT 78.910 -32.970 79.360 -32.860 ;
        RECT 80.760 -32.970 81.210 -32.860 ;
        RECT 82.420 -32.620 82.870 -32.520 ;
        RECT 83.260 -32.620 83.670 -32.190 ;
        RECT 86.420 -32.260 87.970 -32.040 ;
        RECT 88.350 -32.050 88.780 -31.990 ;
        RECT 89.160 -32.040 89.610 -31.990 ;
        RECT 90.210 -32.040 90.710 -31.650 ;
        RECT 89.160 -32.260 90.710 -32.040 ;
        RECT 99.920 -31.650 101.470 -31.430 ;
        RECT 99.920 -32.040 100.420 -31.650 ;
        RECT 101.020 -31.700 101.470 -31.650 ;
        RECT 101.850 -31.700 102.280 -31.640 ;
        RECT 102.660 -31.650 104.210 -31.430 ;
        RECT 106.960 -31.500 107.370 -31.070 ;
        RECT 107.760 -31.170 108.210 -31.070 ;
        RECT 109.420 -30.830 109.870 -30.720 ;
        RECT 111.270 -30.830 111.720 -30.720 ;
        RECT 109.420 -31.070 111.720 -30.830 ;
        RECT 109.420 -31.170 109.870 -31.070 ;
        RECT 110.260 -31.500 110.670 -31.070 ;
        RECT 111.270 -31.140 111.720 -31.070 ;
        RECT 112.670 -30.830 113.120 -30.750 ;
        RECT 113.720 -30.830 114.130 -30.390 ;
        RECT 114.520 -30.830 114.970 -30.720 ;
        RECT 112.670 -31.070 114.970 -30.830 ;
        RECT 112.670 -31.170 113.120 -31.070 ;
        RECT 114.520 -31.170 114.970 -31.070 ;
        RECT 116.160 -30.830 116.610 -30.720 ;
        RECT 117.000 -30.830 117.410 -30.390 ;
        RECT 120.180 -30.660 120.630 -30.380 ;
        RECT 124.000 -30.660 124.450 -30.380 ;
        RECT 133.680 -30.380 135.210 -30.170 ;
        RECT 135.590 -30.260 136.040 -30.170 ;
        RECT 136.420 -30.380 137.950 -30.170 ;
        RECT 118.010 -30.830 118.460 -30.750 ;
        RECT 116.160 -31.070 118.460 -30.830 ;
        RECT 116.160 -31.170 116.610 -31.070 ;
        RECT 118.010 -31.170 118.460 -31.070 ;
        RECT 119.410 -30.830 119.860 -30.720 ;
        RECT 121.260 -30.830 121.710 -30.720 ;
        RECT 119.410 -31.070 121.710 -30.830 ;
        RECT 119.410 -31.140 119.860 -31.070 ;
        RECT 102.660 -31.700 103.110 -31.650 ;
        RECT 101.020 -31.990 103.110 -31.700 ;
        RECT 101.020 -32.040 101.470 -31.990 ;
        RECT 84.270 -32.620 84.720 -32.550 ;
        RECT 82.420 -32.860 84.720 -32.620 ;
        RECT 82.420 -32.970 82.870 -32.860 ;
        RECT 84.270 -32.970 84.720 -32.860 ;
        RECT 85.670 -32.620 86.120 -32.520 ;
        RECT 87.520 -32.620 87.970 -32.520 ;
        RECT 85.670 -32.860 87.970 -32.620 ;
        RECT 85.670 -32.940 86.120 -32.860 ;
        RECT 66.180 -33.520 67.710 -33.310 ;
        RECT 68.090 -33.520 68.540 -33.430 ;
        RECT 68.920 -33.520 70.450 -33.310 ;
        RECT 79.680 -33.310 80.130 -33.030 ;
        RECT 83.500 -33.310 83.950 -33.030 ;
        RECT 86.720 -33.300 87.130 -32.860 ;
        RECT 87.520 -32.970 87.970 -32.860 ;
        RECT 89.160 -32.620 89.610 -32.520 ;
        RECT 91.010 -32.620 91.460 -32.520 ;
        RECT 89.160 -32.860 91.460 -32.620 ;
        RECT 89.160 -32.970 89.610 -32.860 ;
        RECT 90.000 -33.300 90.410 -32.860 ;
        RECT 91.010 -32.940 91.460 -32.860 ;
        RECT 92.410 -32.620 92.860 -32.550 ;
        RECT 93.460 -32.620 93.870 -32.190 ;
        RECT 94.260 -32.620 94.710 -32.520 ;
        RECT 92.410 -32.860 94.710 -32.620 ;
        RECT 92.410 -32.970 92.860 -32.860 ;
        RECT 94.260 -32.970 94.710 -32.860 ;
        RECT 95.920 -32.620 96.370 -32.520 ;
        RECT 96.760 -32.620 97.170 -32.190 ;
        RECT 99.920 -32.260 101.470 -32.040 ;
        RECT 101.850 -32.050 102.280 -31.990 ;
        RECT 102.660 -32.040 103.110 -31.990 ;
        RECT 103.710 -32.040 104.210 -31.650 ;
        RECT 102.660 -32.260 104.210 -32.040 ;
        RECT 113.420 -31.650 114.970 -31.430 ;
        RECT 113.420 -32.040 113.920 -31.650 ;
        RECT 114.520 -31.700 114.970 -31.650 ;
        RECT 115.350 -31.700 115.780 -31.640 ;
        RECT 116.160 -31.650 117.710 -31.430 ;
        RECT 120.460 -31.500 120.870 -31.070 ;
        RECT 121.260 -31.170 121.710 -31.070 ;
        RECT 122.920 -30.830 123.370 -30.720 ;
        RECT 124.770 -30.830 125.220 -30.720 ;
        RECT 122.920 -31.070 125.220 -30.830 ;
        RECT 122.920 -31.170 123.370 -31.070 ;
        RECT 123.760 -31.500 124.170 -31.070 ;
        RECT 124.770 -31.140 125.220 -31.070 ;
        RECT 126.170 -30.830 126.620 -30.750 ;
        RECT 127.220 -30.830 127.630 -30.390 ;
        RECT 128.020 -30.830 128.470 -30.720 ;
        RECT 126.170 -31.070 128.470 -30.830 ;
        RECT 126.170 -31.170 126.620 -31.070 ;
        RECT 128.020 -31.170 128.470 -31.070 ;
        RECT 129.660 -30.830 130.110 -30.720 ;
        RECT 130.500 -30.830 130.910 -30.390 ;
        RECT 133.680 -30.660 134.130 -30.380 ;
        RECT 137.500 -30.660 137.950 -30.380 ;
        RECT 147.180 -30.380 148.710 -30.170 ;
        RECT 149.090 -30.260 149.540 -30.170 ;
        RECT 149.920 -30.380 151.450 -30.170 ;
        RECT 131.510 -30.830 131.960 -30.750 ;
        RECT 129.660 -31.070 131.960 -30.830 ;
        RECT 129.660 -31.170 130.110 -31.070 ;
        RECT 131.510 -31.170 131.960 -31.070 ;
        RECT 132.910 -30.830 133.360 -30.720 ;
        RECT 134.760 -30.830 135.210 -30.720 ;
        RECT 132.910 -31.070 135.210 -30.830 ;
        RECT 132.910 -31.140 133.360 -31.070 ;
        RECT 116.160 -31.700 116.610 -31.650 ;
        RECT 114.520 -31.990 116.610 -31.700 ;
        RECT 114.520 -32.040 114.970 -31.990 ;
        RECT 97.770 -32.620 98.220 -32.550 ;
        RECT 95.920 -32.860 98.220 -32.620 ;
        RECT 95.920 -32.970 96.370 -32.860 ;
        RECT 97.770 -32.970 98.220 -32.860 ;
        RECT 99.170 -32.620 99.620 -32.520 ;
        RECT 101.020 -32.620 101.470 -32.520 ;
        RECT 99.170 -32.860 101.470 -32.620 ;
        RECT 99.170 -32.940 99.620 -32.860 ;
        RECT 79.680 -33.520 81.210 -33.310 ;
        RECT 81.590 -33.520 82.040 -33.430 ;
        RECT 82.420 -33.520 83.950 -33.310 ;
        RECT 93.180 -33.310 93.630 -33.030 ;
        RECT 97.000 -33.310 97.450 -33.030 ;
        RECT 100.220 -33.300 100.630 -32.860 ;
        RECT 101.020 -32.970 101.470 -32.860 ;
        RECT 102.660 -32.620 103.110 -32.520 ;
        RECT 104.510 -32.620 104.960 -32.520 ;
        RECT 102.660 -32.860 104.960 -32.620 ;
        RECT 102.660 -32.970 103.110 -32.860 ;
        RECT 103.500 -33.300 103.910 -32.860 ;
        RECT 104.510 -32.940 104.960 -32.860 ;
        RECT 105.910 -32.620 106.360 -32.550 ;
        RECT 106.960 -32.620 107.370 -32.190 ;
        RECT 107.760 -32.620 108.210 -32.520 ;
        RECT 105.910 -32.860 108.210 -32.620 ;
        RECT 105.910 -32.970 106.360 -32.860 ;
        RECT 107.760 -32.970 108.210 -32.860 ;
        RECT 109.420 -32.620 109.870 -32.520 ;
        RECT 110.260 -32.620 110.670 -32.190 ;
        RECT 113.420 -32.260 114.970 -32.040 ;
        RECT 115.350 -32.050 115.780 -31.990 ;
        RECT 116.160 -32.040 116.610 -31.990 ;
        RECT 117.210 -32.040 117.710 -31.650 ;
        RECT 116.160 -32.260 117.710 -32.040 ;
        RECT 126.920 -31.650 128.470 -31.430 ;
        RECT 126.920 -32.040 127.420 -31.650 ;
        RECT 128.020 -31.700 128.470 -31.650 ;
        RECT 128.850 -31.700 129.280 -31.640 ;
        RECT 129.660 -31.650 131.210 -31.430 ;
        RECT 133.960 -31.500 134.370 -31.070 ;
        RECT 134.760 -31.170 135.210 -31.070 ;
        RECT 136.420 -30.830 136.870 -30.720 ;
        RECT 138.270 -30.830 138.720 -30.720 ;
        RECT 136.420 -31.070 138.720 -30.830 ;
        RECT 136.420 -31.170 136.870 -31.070 ;
        RECT 137.260 -31.500 137.670 -31.070 ;
        RECT 138.270 -31.140 138.720 -31.070 ;
        RECT 139.670 -30.830 140.120 -30.750 ;
        RECT 140.720 -30.830 141.130 -30.390 ;
        RECT 141.520 -30.830 141.970 -30.720 ;
        RECT 139.670 -31.070 141.970 -30.830 ;
        RECT 139.670 -31.170 140.120 -31.070 ;
        RECT 141.520 -31.170 141.970 -31.070 ;
        RECT 143.160 -30.830 143.610 -30.720 ;
        RECT 144.000 -30.830 144.410 -30.390 ;
        RECT 147.180 -30.660 147.630 -30.380 ;
        RECT 151.000 -30.660 151.450 -30.380 ;
        RECT 160.680 -30.380 162.210 -30.170 ;
        RECT 162.590 -30.260 163.040 -30.170 ;
        RECT 163.420 -30.380 164.950 -30.170 ;
        RECT 145.010 -30.830 145.460 -30.750 ;
        RECT 143.160 -31.070 145.460 -30.830 ;
        RECT 143.160 -31.170 143.610 -31.070 ;
        RECT 145.010 -31.170 145.460 -31.070 ;
        RECT 146.410 -30.830 146.860 -30.720 ;
        RECT 148.260 -30.830 148.710 -30.720 ;
        RECT 146.410 -31.070 148.710 -30.830 ;
        RECT 146.410 -31.140 146.860 -31.070 ;
        RECT 129.660 -31.700 130.110 -31.650 ;
        RECT 128.020 -31.990 130.110 -31.700 ;
        RECT 128.020 -32.040 128.470 -31.990 ;
        RECT 111.270 -32.620 111.720 -32.550 ;
        RECT 109.420 -32.860 111.720 -32.620 ;
        RECT 109.420 -32.970 109.870 -32.860 ;
        RECT 111.270 -32.970 111.720 -32.860 ;
        RECT 112.670 -32.620 113.120 -32.520 ;
        RECT 114.520 -32.620 114.970 -32.520 ;
        RECT 112.670 -32.860 114.970 -32.620 ;
        RECT 112.670 -32.940 113.120 -32.860 ;
        RECT 93.180 -33.520 94.710 -33.310 ;
        RECT 95.090 -33.520 95.540 -33.430 ;
        RECT 95.920 -33.520 97.450 -33.310 ;
        RECT 106.680 -33.310 107.130 -33.030 ;
        RECT 110.500 -33.310 110.950 -33.030 ;
        RECT 113.720 -33.300 114.130 -32.860 ;
        RECT 114.520 -32.970 114.970 -32.860 ;
        RECT 116.160 -32.620 116.610 -32.520 ;
        RECT 118.010 -32.620 118.460 -32.520 ;
        RECT 116.160 -32.860 118.460 -32.620 ;
        RECT 116.160 -32.970 116.610 -32.860 ;
        RECT 117.000 -33.300 117.410 -32.860 ;
        RECT 118.010 -32.940 118.460 -32.860 ;
        RECT 119.410 -32.620 119.860 -32.550 ;
        RECT 120.460 -32.620 120.870 -32.190 ;
        RECT 121.260 -32.620 121.710 -32.520 ;
        RECT 119.410 -32.860 121.710 -32.620 ;
        RECT 119.410 -32.970 119.860 -32.860 ;
        RECT 121.260 -32.970 121.710 -32.860 ;
        RECT 122.920 -32.620 123.370 -32.520 ;
        RECT 123.760 -32.620 124.170 -32.190 ;
        RECT 126.920 -32.260 128.470 -32.040 ;
        RECT 128.850 -32.050 129.280 -31.990 ;
        RECT 129.660 -32.040 130.110 -31.990 ;
        RECT 130.710 -32.040 131.210 -31.650 ;
        RECT 129.660 -32.260 131.210 -32.040 ;
        RECT 140.420 -31.650 141.970 -31.430 ;
        RECT 140.420 -32.040 140.920 -31.650 ;
        RECT 141.520 -31.700 141.970 -31.650 ;
        RECT 142.350 -31.700 142.780 -31.640 ;
        RECT 143.160 -31.650 144.710 -31.430 ;
        RECT 147.460 -31.500 147.870 -31.070 ;
        RECT 148.260 -31.170 148.710 -31.070 ;
        RECT 149.920 -30.830 150.370 -30.720 ;
        RECT 151.770 -30.830 152.220 -30.720 ;
        RECT 149.920 -31.070 152.220 -30.830 ;
        RECT 149.920 -31.170 150.370 -31.070 ;
        RECT 150.760 -31.500 151.170 -31.070 ;
        RECT 151.770 -31.140 152.220 -31.070 ;
        RECT 153.170 -30.830 153.620 -30.750 ;
        RECT 154.220 -30.830 154.630 -30.390 ;
        RECT 155.020 -30.830 155.470 -30.720 ;
        RECT 153.170 -31.070 155.470 -30.830 ;
        RECT 153.170 -31.170 153.620 -31.070 ;
        RECT 155.020 -31.170 155.470 -31.070 ;
        RECT 156.660 -30.830 157.110 -30.720 ;
        RECT 157.500 -30.830 157.910 -30.390 ;
        RECT 160.680 -30.660 161.130 -30.380 ;
        RECT 164.500 -30.660 164.950 -30.380 ;
        RECT 174.180 -30.380 175.710 -30.170 ;
        RECT 176.090 -30.260 176.540 -30.170 ;
        RECT 176.920 -30.380 178.450 -30.170 ;
        RECT 158.510 -30.830 158.960 -30.750 ;
        RECT 156.660 -31.070 158.960 -30.830 ;
        RECT 156.660 -31.170 157.110 -31.070 ;
        RECT 158.510 -31.170 158.960 -31.070 ;
        RECT 159.910 -30.830 160.360 -30.720 ;
        RECT 161.760 -30.830 162.210 -30.720 ;
        RECT 159.910 -31.070 162.210 -30.830 ;
        RECT 159.910 -31.140 160.360 -31.070 ;
        RECT 143.160 -31.700 143.610 -31.650 ;
        RECT 141.520 -31.990 143.610 -31.700 ;
        RECT 141.520 -32.040 141.970 -31.990 ;
        RECT 124.770 -32.620 125.220 -32.550 ;
        RECT 122.920 -32.860 125.220 -32.620 ;
        RECT 122.920 -32.970 123.370 -32.860 ;
        RECT 124.770 -32.970 125.220 -32.860 ;
        RECT 126.170 -32.620 126.620 -32.520 ;
        RECT 128.020 -32.620 128.470 -32.520 ;
        RECT 126.170 -32.860 128.470 -32.620 ;
        RECT 126.170 -32.940 126.620 -32.860 ;
        RECT 106.680 -33.520 108.210 -33.310 ;
        RECT 108.590 -33.520 109.040 -33.430 ;
        RECT 109.420 -33.520 110.950 -33.310 ;
        RECT 120.180 -33.310 120.630 -33.030 ;
        RECT 124.000 -33.310 124.450 -33.030 ;
        RECT 127.220 -33.300 127.630 -32.860 ;
        RECT 128.020 -32.970 128.470 -32.860 ;
        RECT 129.660 -32.620 130.110 -32.520 ;
        RECT 131.510 -32.620 131.960 -32.520 ;
        RECT 129.660 -32.860 131.960 -32.620 ;
        RECT 129.660 -32.970 130.110 -32.860 ;
        RECT 130.500 -33.300 130.910 -32.860 ;
        RECT 131.510 -32.940 131.960 -32.860 ;
        RECT 132.910 -32.620 133.360 -32.550 ;
        RECT 133.960 -32.620 134.370 -32.190 ;
        RECT 134.760 -32.620 135.210 -32.520 ;
        RECT 132.910 -32.860 135.210 -32.620 ;
        RECT 132.910 -32.970 133.360 -32.860 ;
        RECT 134.760 -32.970 135.210 -32.860 ;
        RECT 136.420 -32.620 136.870 -32.520 ;
        RECT 137.260 -32.620 137.670 -32.190 ;
        RECT 140.420 -32.260 141.970 -32.040 ;
        RECT 142.350 -32.050 142.780 -31.990 ;
        RECT 143.160 -32.040 143.610 -31.990 ;
        RECT 144.210 -32.040 144.710 -31.650 ;
        RECT 143.160 -32.260 144.710 -32.040 ;
        RECT 153.920 -31.650 155.470 -31.430 ;
        RECT 153.920 -32.040 154.420 -31.650 ;
        RECT 155.020 -31.700 155.470 -31.650 ;
        RECT 155.850 -31.700 156.280 -31.640 ;
        RECT 156.660 -31.650 158.210 -31.430 ;
        RECT 160.960 -31.500 161.370 -31.070 ;
        RECT 161.760 -31.170 162.210 -31.070 ;
        RECT 163.420 -30.830 163.870 -30.720 ;
        RECT 165.270 -30.830 165.720 -30.720 ;
        RECT 163.420 -31.070 165.720 -30.830 ;
        RECT 163.420 -31.170 163.870 -31.070 ;
        RECT 164.260 -31.500 164.670 -31.070 ;
        RECT 165.270 -31.140 165.720 -31.070 ;
        RECT 166.670 -30.830 167.120 -30.750 ;
        RECT 167.720 -30.830 168.130 -30.390 ;
        RECT 168.520 -30.830 168.970 -30.720 ;
        RECT 166.670 -31.070 168.970 -30.830 ;
        RECT 166.670 -31.170 167.120 -31.070 ;
        RECT 168.520 -31.170 168.970 -31.070 ;
        RECT 170.160 -30.830 170.610 -30.720 ;
        RECT 171.000 -30.830 171.410 -30.390 ;
        RECT 174.180 -30.660 174.630 -30.380 ;
        RECT 178.000 -30.660 178.450 -30.380 ;
        RECT 187.680 -30.380 189.210 -30.170 ;
        RECT 189.590 -30.260 190.040 -30.170 ;
        RECT 190.420 -30.380 191.950 -30.170 ;
        RECT 172.010 -30.830 172.460 -30.750 ;
        RECT 170.160 -31.070 172.460 -30.830 ;
        RECT 170.160 -31.170 170.610 -31.070 ;
        RECT 172.010 -31.170 172.460 -31.070 ;
        RECT 173.410 -30.830 173.860 -30.720 ;
        RECT 175.260 -30.830 175.710 -30.720 ;
        RECT 173.410 -31.070 175.710 -30.830 ;
        RECT 173.410 -31.140 173.860 -31.070 ;
        RECT 156.660 -31.700 157.110 -31.650 ;
        RECT 155.020 -31.990 157.110 -31.700 ;
        RECT 155.020 -32.040 155.470 -31.990 ;
        RECT 138.270 -32.620 138.720 -32.550 ;
        RECT 136.420 -32.860 138.720 -32.620 ;
        RECT 136.420 -32.970 136.870 -32.860 ;
        RECT 138.270 -32.970 138.720 -32.860 ;
        RECT 139.670 -32.620 140.120 -32.520 ;
        RECT 141.520 -32.620 141.970 -32.520 ;
        RECT 139.670 -32.860 141.970 -32.620 ;
        RECT 139.670 -32.940 140.120 -32.860 ;
        RECT 120.180 -33.520 121.710 -33.310 ;
        RECT 122.090 -33.520 122.540 -33.430 ;
        RECT 122.920 -33.520 124.450 -33.310 ;
        RECT 133.680 -33.310 134.130 -33.030 ;
        RECT 137.500 -33.310 137.950 -33.030 ;
        RECT 140.720 -33.300 141.130 -32.860 ;
        RECT 141.520 -32.970 141.970 -32.860 ;
        RECT 143.160 -32.620 143.610 -32.520 ;
        RECT 145.010 -32.620 145.460 -32.520 ;
        RECT 143.160 -32.860 145.460 -32.620 ;
        RECT 143.160 -32.970 143.610 -32.860 ;
        RECT 144.000 -33.300 144.410 -32.860 ;
        RECT 145.010 -32.940 145.460 -32.860 ;
        RECT 146.410 -32.620 146.860 -32.550 ;
        RECT 147.460 -32.620 147.870 -32.190 ;
        RECT 148.260 -32.620 148.710 -32.520 ;
        RECT 146.410 -32.860 148.710 -32.620 ;
        RECT 146.410 -32.970 146.860 -32.860 ;
        RECT 148.260 -32.970 148.710 -32.860 ;
        RECT 149.920 -32.620 150.370 -32.520 ;
        RECT 150.760 -32.620 151.170 -32.190 ;
        RECT 153.920 -32.260 155.470 -32.040 ;
        RECT 155.850 -32.050 156.280 -31.990 ;
        RECT 156.660 -32.040 157.110 -31.990 ;
        RECT 157.710 -32.040 158.210 -31.650 ;
        RECT 156.660 -32.260 158.210 -32.040 ;
        RECT 167.420 -31.650 168.970 -31.430 ;
        RECT 167.420 -32.040 167.920 -31.650 ;
        RECT 168.520 -31.700 168.970 -31.650 ;
        RECT 169.350 -31.700 169.780 -31.640 ;
        RECT 170.160 -31.650 171.710 -31.430 ;
        RECT 174.460 -31.500 174.870 -31.070 ;
        RECT 175.260 -31.170 175.710 -31.070 ;
        RECT 176.920 -30.830 177.370 -30.720 ;
        RECT 178.770 -30.830 179.220 -30.720 ;
        RECT 176.920 -31.070 179.220 -30.830 ;
        RECT 176.920 -31.170 177.370 -31.070 ;
        RECT 177.760 -31.500 178.170 -31.070 ;
        RECT 178.770 -31.140 179.220 -31.070 ;
        RECT 180.170 -30.830 180.620 -30.750 ;
        RECT 181.220 -30.830 181.630 -30.390 ;
        RECT 182.020 -30.830 182.470 -30.720 ;
        RECT 180.170 -31.070 182.470 -30.830 ;
        RECT 180.170 -31.170 180.620 -31.070 ;
        RECT 182.020 -31.170 182.470 -31.070 ;
        RECT 183.660 -30.830 184.110 -30.720 ;
        RECT 184.500 -30.830 184.910 -30.390 ;
        RECT 187.680 -30.660 188.130 -30.380 ;
        RECT 191.500 -30.660 191.950 -30.380 ;
        RECT 201.180 -30.380 202.710 -30.170 ;
        RECT 203.090 -30.260 203.540 -30.170 ;
        RECT 203.920 -30.380 205.450 -30.170 ;
        RECT 185.510 -30.830 185.960 -30.750 ;
        RECT 183.660 -31.070 185.960 -30.830 ;
        RECT 183.660 -31.170 184.110 -31.070 ;
        RECT 185.510 -31.170 185.960 -31.070 ;
        RECT 186.910 -30.830 187.360 -30.720 ;
        RECT 188.760 -30.830 189.210 -30.720 ;
        RECT 186.910 -31.070 189.210 -30.830 ;
        RECT 186.910 -31.140 187.360 -31.070 ;
        RECT 170.160 -31.700 170.610 -31.650 ;
        RECT 168.520 -31.990 170.610 -31.700 ;
        RECT 168.520 -32.040 168.970 -31.990 ;
        RECT 151.770 -32.620 152.220 -32.550 ;
        RECT 149.920 -32.860 152.220 -32.620 ;
        RECT 149.920 -32.970 150.370 -32.860 ;
        RECT 151.770 -32.970 152.220 -32.860 ;
        RECT 153.170 -32.620 153.620 -32.520 ;
        RECT 155.020 -32.620 155.470 -32.520 ;
        RECT 153.170 -32.860 155.470 -32.620 ;
        RECT 153.170 -32.940 153.620 -32.860 ;
        RECT 133.680 -33.520 135.210 -33.310 ;
        RECT 135.590 -33.520 136.040 -33.430 ;
        RECT 136.420 -33.520 137.950 -33.310 ;
        RECT 147.180 -33.310 147.630 -33.030 ;
        RECT 151.000 -33.310 151.450 -33.030 ;
        RECT 154.220 -33.300 154.630 -32.860 ;
        RECT 155.020 -32.970 155.470 -32.860 ;
        RECT 156.660 -32.620 157.110 -32.520 ;
        RECT 158.510 -32.620 158.960 -32.520 ;
        RECT 156.660 -32.860 158.960 -32.620 ;
        RECT 156.660 -32.970 157.110 -32.860 ;
        RECT 157.500 -33.300 157.910 -32.860 ;
        RECT 158.510 -32.940 158.960 -32.860 ;
        RECT 159.910 -32.620 160.360 -32.550 ;
        RECT 160.960 -32.620 161.370 -32.190 ;
        RECT 161.760 -32.620 162.210 -32.520 ;
        RECT 159.910 -32.860 162.210 -32.620 ;
        RECT 159.910 -32.970 160.360 -32.860 ;
        RECT 161.760 -32.970 162.210 -32.860 ;
        RECT 163.420 -32.620 163.870 -32.520 ;
        RECT 164.260 -32.620 164.670 -32.190 ;
        RECT 167.420 -32.260 168.970 -32.040 ;
        RECT 169.350 -32.050 169.780 -31.990 ;
        RECT 170.160 -32.040 170.610 -31.990 ;
        RECT 171.210 -32.040 171.710 -31.650 ;
        RECT 170.160 -32.260 171.710 -32.040 ;
        RECT 180.920 -31.650 182.470 -31.430 ;
        RECT 180.920 -32.040 181.420 -31.650 ;
        RECT 182.020 -31.700 182.470 -31.650 ;
        RECT 182.850 -31.700 183.280 -31.640 ;
        RECT 183.660 -31.650 185.210 -31.430 ;
        RECT 187.960 -31.500 188.370 -31.070 ;
        RECT 188.760 -31.170 189.210 -31.070 ;
        RECT 190.420 -30.830 190.870 -30.720 ;
        RECT 192.270 -30.830 192.720 -30.720 ;
        RECT 190.420 -31.070 192.720 -30.830 ;
        RECT 190.420 -31.170 190.870 -31.070 ;
        RECT 191.260 -31.500 191.670 -31.070 ;
        RECT 192.270 -31.140 192.720 -31.070 ;
        RECT 193.670 -30.830 194.120 -30.750 ;
        RECT 194.720 -30.830 195.130 -30.390 ;
        RECT 195.520 -30.830 195.970 -30.720 ;
        RECT 193.670 -31.070 195.970 -30.830 ;
        RECT 193.670 -31.170 194.120 -31.070 ;
        RECT 195.520 -31.170 195.970 -31.070 ;
        RECT 197.160 -30.830 197.610 -30.720 ;
        RECT 198.000 -30.830 198.410 -30.390 ;
        RECT 201.180 -30.660 201.630 -30.380 ;
        RECT 205.000 -30.660 205.450 -30.380 ;
        RECT 214.680 -30.380 216.210 -30.170 ;
        RECT 216.590 -30.260 217.030 -30.170 ;
        RECT 199.010 -30.830 199.460 -30.750 ;
        RECT 197.160 -31.070 199.460 -30.830 ;
        RECT 197.160 -31.170 197.610 -31.070 ;
        RECT 199.010 -31.170 199.460 -31.070 ;
        RECT 200.410 -30.830 200.860 -30.720 ;
        RECT 202.260 -30.830 202.710 -30.720 ;
        RECT 200.410 -31.070 202.710 -30.830 ;
        RECT 200.410 -31.140 200.860 -31.070 ;
        RECT 183.660 -31.700 184.110 -31.650 ;
        RECT 182.020 -31.990 184.110 -31.700 ;
        RECT 182.020 -32.040 182.470 -31.990 ;
        RECT 165.270 -32.620 165.720 -32.550 ;
        RECT 163.420 -32.860 165.720 -32.620 ;
        RECT 163.420 -32.970 163.870 -32.860 ;
        RECT 165.270 -32.970 165.720 -32.860 ;
        RECT 166.670 -32.620 167.120 -32.520 ;
        RECT 168.520 -32.620 168.970 -32.520 ;
        RECT 166.670 -32.860 168.970 -32.620 ;
        RECT 166.670 -32.940 167.120 -32.860 ;
        RECT 147.180 -33.520 148.710 -33.310 ;
        RECT 149.090 -33.520 149.540 -33.430 ;
        RECT 149.920 -33.520 151.450 -33.310 ;
        RECT 160.680 -33.310 161.130 -33.030 ;
        RECT 164.500 -33.310 164.950 -33.030 ;
        RECT 167.720 -33.300 168.130 -32.860 ;
        RECT 168.520 -32.970 168.970 -32.860 ;
        RECT 170.160 -32.620 170.610 -32.520 ;
        RECT 172.010 -32.620 172.460 -32.520 ;
        RECT 170.160 -32.860 172.460 -32.620 ;
        RECT 170.160 -32.970 170.610 -32.860 ;
        RECT 171.000 -33.300 171.410 -32.860 ;
        RECT 172.010 -32.940 172.460 -32.860 ;
        RECT 173.410 -32.620 173.860 -32.550 ;
        RECT 174.460 -32.620 174.870 -32.190 ;
        RECT 175.260 -32.620 175.710 -32.520 ;
        RECT 173.410 -32.860 175.710 -32.620 ;
        RECT 173.410 -32.970 173.860 -32.860 ;
        RECT 175.260 -32.970 175.710 -32.860 ;
        RECT 176.920 -32.620 177.370 -32.520 ;
        RECT 177.760 -32.620 178.170 -32.190 ;
        RECT 180.920 -32.260 182.470 -32.040 ;
        RECT 182.850 -32.050 183.280 -31.990 ;
        RECT 183.660 -32.040 184.110 -31.990 ;
        RECT 184.710 -32.040 185.210 -31.650 ;
        RECT 183.660 -32.260 185.210 -32.040 ;
        RECT 194.420 -31.650 195.970 -31.430 ;
        RECT 194.420 -32.040 194.920 -31.650 ;
        RECT 195.520 -31.700 195.970 -31.650 ;
        RECT 196.350 -31.700 196.780 -31.640 ;
        RECT 197.160 -31.650 198.710 -31.430 ;
        RECT 201.460 -31.500 201.870 -31.070 ;
        RECT 202.260 -31.170 202.710 -31.070 ;
        RECT 203.920 -30.830 204.370 -30.720 ;
        RECT 205.770 -30.830 206.220 -30.720 ;
        RECT 203.920 -31.070 206.220 -30.830 ;
        RECT 203.920 -31.170 204.370 -31.070 ;
        RECT 204.760 -31.500 205.170 -31.070 ;
        RECT 205.770 -31.140 206.220 -31.070 ;
        RECT 207.170 -30.830 207.620 -30.750 ;
        RECT 208.220 -30.830 208.630 -30.390 ;
        RECT 209.020 -30.830 209.470 -30.720 ;
        RECT 207.170 -31.070 209.470 -30.830 ;
        RECT 207.170 -31.170 207.620 -31.070 ;
        RECT 209.020 -31.170 209.470 -31.070 ;
        RECT 210.660 -30.830 211.110 -30.720 ;
        RECT 211.500 -30.830 211.910 -30.390 ;
        RECT 214.680 -30.660 215.130 -30.380 ;
        RECT 212.510 -30.830 212.960 -30.750 ;
        RECT 210.660 -31.070 212.960 -30.830 ;
        RECT 210.660 -31.170 211.110 -31.070 ;
        RECT 212.510 -31.170 212.960 -31.070 ;
        RECT 213.910 -30.830 214.360 -30.720 ;
        RECT 215.760 -30.830 216.210 -30.720 ;
        RECT 213.910 -31.070 216.210 -30.830 ;
        RECT 213.910 -31.140 214.360 -31.070 ;
        RECT 197.160 -31.700 197.610 -31.650 ;
        RECT 195.520 -31.990 197.610 -31.700 ;
        RECT 195.520 -32.040 195.970 -31.990 ;
        RECT 178.770 -32.620 179.220 -32.550 ;
        RECT 176.920 -32.860 179.220 -32.620 ;
        RECT 176.920 -32.970 177.370 -32.860 ;
        RECT 178.770 -32.970 179.220 -32.860 ;
        RECT 180.170 -32.620 180.620 -32.520 ;
        RECT 182.020 -32.620 182.470 -32.520 ;
        RECT 180.170 -32.860 182.470 -32.620 ;
        RECT 180.170 -32.940 180.620 -32.860 ;
        RECT 160.680 -33.520 162.210 -33.310 ;
        RECT 162.590 -33.520 163.040 -33.430 ;
        RECT 163.420 -33.520 164.950 -33.310 ;
        RECT 174.180 -33.310 174.630 -33.030 ;
        RECT 178.000 -33.310 178.450 -33.030 ;
        RECT 181.220 -33.300 181.630 -32.860 ;
        RECT 182.020 -32.970 182.470 -32.860 ;
        RECT 183.660 -32.620 184.110 -32.520 ;
        RECT 185.510 -32.620 185.960 -32.520 ;
        RECT 183.660 -32.860 185.960 -32.620 ;
        RECT 183.660 -32.970 184.110 -32.860 ;
        RECT 184.500 -33.300 184.910 -32.860 ;
        RECT 185.510 -32.940 185.960 -32.860 ;
        RECT 186.910 -32.620 187.360 -32.550 ;
        RECT 187.960 -32.620 188.370 -32.190 ;
        RECT 188.760 -32.620 189.210 -32.520 ;
        RECT 186.910 -32.860 189.210 -32.620 ;
        RECT 186.910 -32.970 187.360 -32.860 ;
        RECT 188.760 -32.970 189.210 -32.860 ;
        RECT 190.420 -32.620 190.870 -32.520 ;
        RECT 191.260 -32.620 191.670 -32.190 ;
        RECT 194.420 -32.260 195.970 -32.040 ;
        RECT 196.350 -32.050 196.780 -31.990 ;
        RECT 197.160 -32.040 197.610 -31.990 ;
        RECT 198.210 -32.040 198.710 -31.650 ;
        RECT 197.160 -32.260 198.710 -32.040 ;
        RECT 207.920 -31.650 209.470 -31.430 ;
        RECT 207.920 -32.040 208.420 -31.650 ;
        RECT 209.020 -31.700 209.470 -31.650 ;
        RECT 209.850 -31.700 210.280 -31.640 ;
        RECT 210.660 -31.650 212.210 -31.430 ;
        RECT 214.960 -31.500 215.370 -31.070 ;
        RECT 215.760 -31.170 216.210 -31.070 ;
        RECT 210.660 -31.700 211.110 -31.650 ;
        RECT 209.020 -31.990 211.110 -31.700 ;
        RECT 209.020 -32.040 209.470 -31.990 ;
        RECT 192.270 -32.620 192.720 -32.550 ;
        RECT 190.420 -32.860 192.720 -32.620 ;
        RECT 190.420 -32.970 190.870 -32.860 ;
        RECT 192.270 -32.970 192.720 -32.860 ;
        RECT 193.670 -32.620 194.120 -32.520 ;
        RECT 195.520 -32.620 195.970 -32.520 ;
        RECT 193.670 -32.860 195.970 -32.620 ;
        RECT 193.670 -32.940 194.120 -32.860 ;
        RECT 174.180 -33.520 175.710 -33.310 ;
        RECT 176.090 -33.520 176.540 -33.430 ;
        RECT 176.920 -33.520 178.450 -33.310 ;
        RECT 187.680 -33.310 188.130 -33.030 ;
        RECT 191.500 -33.310 191.950 -33.030 ;
        RECT 194.720 -33.300 195.130 -32.860 ;
        RECT 195.520 -32.970 195.970 -32.860 ;
        RECT 197.160 -32.620 197.610 -32.520 ;
        RECT 199.010 -32.620 199.460 -32.520 ;
        RECT 197.160 -32.860 199.460 -32.620 ;
        RECT 197.160 -32.970 197.610 -32.860 ;
        RECT 198.000 -33.300 198.410 -32.860 ;
        RECT 199.010 -32.940 199.460 -32.860 ;
        RECT 200.410 -32.620 200.860 -32.550 ;
        RECT 201.460 -32.620 201.870 -32.190 ;
        RECT 202.260 -32.620 202.710 -32.520 ;
        RECT 200.410 -32.860 202.710 -32.620 ;
        RECT 200.410 -32.970 200.860 -32.860 ;
        RECT 202.260 -32.970 202.710 -32.860 ;
        RECT 203.920 -32.620 204.370 -32.520 ;
        RECT 204.760 -32.620 205.170 -32.190 ;
        RECT 207.920 -32.260 209.470 -32.040 ;
        RECT 209.850 -32.050 210.280 -31.990 ;
        RECT 210.660 -32.040 211.110 -31.990 ;
        RECT 211.710 -32.040 212.210 -31.650 ;
        RECT 210.660 -32.260 212.210 -32.040 ;
        RECT 205.770 -32.620 206.220 -32.550 ;
        RECT 203.920 -32.860 206.220 -32.620 ;
        RECT 203.920 -32.970 204.370 -32.860 ;
        RECT 205.770 -32.970 206.220 -32.860 ;
        RECT 207.170 -32.620 207.620 -32.520 ;
        RECT 209.020 -32.620 209.470 -32.520 ;
        RECT 207.170 -32.860 209.470 -32.620 ;
        RECT 207.170 -32.940 207.620 -32.860 ;
        RECT 187.680 -33.520 189.210 -33.310 ;
        RECT 189.590 -33.520 190.040 -33.430 ;
        RECT 190.420 -33.520 191.950 -33.310 ;
        RECT 201.180 -33.310 201.630 -33.030 ;
        RECT 205.000 -33.310 205.450 -33.030 ;
        RECT 208.220 -33.300 208.630 -32.860 ;
        RECT 209.020 -32.970 209.470 -32.860 ;
        RECT 210.660 -32.620 211.110 -32.520 ;
        RECT 212.510 -32.620 212.960 -32.520 ;
        RECT 210.660 -32.860 212.960 -32.620 ;
        RECT 210.660 -32.970 211.110 -32.860 ;
        RECT 211.500 -33.300 211.910 -32.860 ;
        RECT 212.510 -32.940 212.960 -32.860 ;
        RECT 213.910 -32.620 214.360 -32.550 ;
        RECT 214.960 -32.620 215.370 -32.190 ;
        RECT 215.760 -32.620 216.210 -32.520 ;
        RECT 213.910 -32.860 216.210 -32.620 ;
        RECT 213.910 -32.970 214.360 -32.860 ;
        RECT 215.760 -32.970 216.210 -32.860 ;
        RECT 201.180 -33.520 202.710 -33.310 ;
        RECT 203.090 -33.520 203.540 -33.430 ;
        RECT 203.920 -33.520 205.450 -33.310 ;
        RECT 214.680 -33.310 215.130 -33.030 ;
        RECT 214.680 -33.520 216.210 -33.310 ;
        RECT 216.590 -33.520 217.030 -33.430 ;
        RECT 13.260 -33.780 15.370 -33.520 ;
        RECT 26.760 -33.780 28.870 -33.520 ;
        RECT 40.260 -33.780 42.370 -33.520 ;
        RECT 53.760 -33.780 55.870 -33.520 ;
        RECT 67.260 -33.780 69.370 -33.520 ;
        RECT 80.760 -33.780 82.870 -33.520 ;
        RECT 94.260 -33.780 96.370 -33.520 ;
        RECT 107.760 -33.780 109.870 -33.520 ;
        RECT 121.260 -33.780 123.370 -33.520 ;
        RECT 134.760 -33.780 136.870 -33.520 ;
        RECT 148.260 -33.780 150.370 -33.520 ;
        RECT 161.760 -33.780 163.870 -33.520 ;
        RECT 175.260 -33.780 177.370 -33.520 ;
        RECT 188.760 -33.780 190.870 -33.520 ;
        RECT 202.260 -33.780 204.370 -33.520 ;
        RECT 215.760 -33.780 217.030 -33.520 ;
        RECT 12.180 -33.990 13.710 -33.780 ;
        RECT 14.090 -33.870 14.540 -33.780 ;
        RECT 14.920 -33.990 16.450 -33.780 ;
        RECT 1.420 -34.440 1.870 -34.330 ;
        RECT 3.270 -34.440 3.720 -34.330 ;
        RECT 1.420 -34.680 3.720 -34.440 ;
        RECT 1.420 -34.780 1.870 -34.680 ;
        RECT 2.260 -35.110 2.670 -34.680 ;
        RECT 3.270 -34.750 3.720 -34.680 ;
        RECT 4.670 -34.440 5.120 -34.360 ;
        RECT 5.720 -34.440 6.130 -34.000 ;
        RECT 6.520 -34.440 6.970 -34.330 ;
        RECT 4.670 -34.680 6.970 -34.440 ;
        RECT 4.670 -34.780 5.120 -34.680 ;
        RECT 6.520 -34.780 6.970 -34.680 ;
        RECT 8.160 -34.440 8.610 -34.330 ;
        RECT 9.000 -34.440 9.410 -34.000 ;
        RECT 12.180 -34.270 12.630 -33.990 ;
        RECT 16.000 -34.270 16.450 -33.990 ;
        RECT 25.680 -33.990 27.210 -33.780 ;
        RECT 27.590 -33.870 28.040 -33.780 ;
        RECT 28.420 -33.990 29.950 -33.780 ;
        RECT 10.010 -34.440 10.460 -34.360 ;
        RECT 8.160 -34.680 10.460 -34.440 ;
        RECT 8.160 -34.780 8.610 -34.680 ;
        RECT 10.010 -34.780 10.460 -34.680 ;
        RECT 11.410 -34.440 11.860 -34.330 ;
        RECT 13.260 -34.440 13.710 -34.330 ;
        RECT 11.410 -34.680 13.710 -34.440 ;
        RECT 11.410 -34.750 11.860 -34.680 ;
        RECT 5.420 -35.260 6.970 -35.040 ;
        RECT 5.420 -35.650 5.920 -35.260 ;
        RECT 6.520 -35.310 6.970 -35.260 ;
        RECT 7.350 -35.310 7.780 -35.250 ;
        RECT 8.160 -35.260 9.710 -35.040 ;
        RECT 12.460 -35.110 12.870 -34.680 ;
        RECT 13.260 -34.780 13.710 -34.680 ;
        RECT 14.920 -34.440 15.370 -34.330 ;
        RECT 16.770 -34.440 17.220 -34.330 ;
        RECT 14.920 -34.680 17.220 -34.440 ;
        RECT 14.920 -34.780 15.370 -34.680 ;
        RECT 15.760 -35.110 16.170 -34.680 ;
        RECT 16.770 -34.750 17.220 -34.680 ;
        RECT 18.170 -34.440 18.620 -34.360 ;
        RECT 19.220 -34.440 19.630 -34.000 ;
        RECT 20.020 -34.440 20.470 -34.330 ;
        RECT 18.170 -34.680 20.470 -34.440 ;
        RECT 18.170 -34.780 18.620 -34.680 ;
        RECT 20.020 -34.780 20.470 -34.680 ;
        RECT 21.660 -34.440 22.110 -34.330 ;
        RECT 22.500 -34.440 22.910 -34.000 ;
        RECT 25.680 -34.270 26.130 -33.990 ;
        RECT 29.500 -34.270 29.950 -33.990 ;
        RECT 39.180 -33.990 40.710 -33.780 ;
        RECT 41.090 -33.870 41.540 -33.780 ;
        RECT 41.920 -33.990 43.450 -33.780 ;
        RECT 23.510 -34.440 23.960 -34.360 ;
        RECT 21.660 -34.680 23.960 -34.440 ;
        RECT 21.660 -34.780 22.110 -34.680 ;
        RECT 23.510 -34.780 23.960 -34.680 ;
        RECT 24.910 -34.440 25.360 -34.330 ;
        RECT 26.760 -34.440 27.210 -34.330 ;
        RECT 24.910 -34.680 27.210 -34.440 ;
        RECT 24.910 -34.750 25.360 -34.680 ;
        RECT 8.160 -35.310 8.610 -35.260 ;
        RECT 6.520 -35.600 8.610 -35.310 ;
        RECT 6.520 -35.650 6.970 -35.600 ;
        RECT 1.420 -36.230 1.870 -36.130 ;
        RECT 2.260 -36.230 2.670 -35.800 ;
        RECT 5.420 -35.870 6.970 -35.650 ;
        RECT 7.350 -35.660 7.780 -35.600 ;
        RECT 8.160 -35.650 8.610 -35.600 ;
        RECT 9.210 -35.650 9.710 -35.260 ;
        RECT 8.160 -35.870 9.710 -35.650 ;
        RECT 18.920 -35.260 20.470 -35.040 ;
        RECT 18.920 -35.650 19.420 -35.260 ;
        RECT 20.020 -35.310 20.470 -35.260 ;
        RECT 20.850 -35.310 21.280 -35.250 ;
        RECT 21.660 -35.260 23.210 -35.040 ;
        RECT 25.960 -35.110 26.370 -34.680 ;
        RECT 26.760 -34.780 27.210 -34.680 ;
        RECT 28.420 -34.440 28.870 -34.330 ;
        RECT 30.270 -34.440 30.720 -34.330 ;
        RECT 28.420 -34.680 30.720 -34.440 ;
        RECT 28.420 -34.780 28.870 -34.680 ;
        RECT 29.260 -35.110 29.670 -34.680 ;
        RECT 30.270 -34.750 30.720 -34.680 ;
        RECT 31.670 -34.440 32.120 -34.360 ;
        RECT 32.720 -34.440 33.130 -34.000 ;
        RECT 33.520 -34.440 33.970 -34.330 ;
        RECT 31.670 -34.680 33.970 -34.440 ;
        RECT 31.670 -34.780 32.120 -34.680 ;
        RECT 33.520 -34.780 33.970 -34.680 ;
        RECT 35.160 -34.440 35.610 -34.330 ;
        RECT 36.000 -34.440 36.410 -34.000 ;
        RECT 39.180 -34.270 39.630 -33.990 ;
        RECT 43.000 -34.270 43.450 -33.990 ;
        RECT 52.680 -33.990 54.210 -33.780 ;
        RECT 54.590 -33.870 55.040 -33.780 ;
        RECT 55.420 -33.990 56.950 -33.780 ;
        RECT 37.010 -34.440 37.460 -34.360 ;
        RECT 35.160 -34.680 37.460 -34.440 ;
        RECT 35.160 -34.780 35.610 -34.680 ;
        RECT 37.010 -34.780 37.460 -34.680 ;
        RECT 38.410 -34.440 38.860 -34.330 ;
        RECT 40.260 -34.440 40.710 -34.330 ;
        RECT 38.410 -34.680 40.710 -34.440 ;
        RECT 38.410 -34.750 38.860 -34.680 ;
        RECT 21.660 -35.310 22.110 -35.260 ;
        RECT 20.020 -35.600 22.110 -35.310 ;
        RECT 20.020 -35.650 20.470 -35.600 ;
        RECT 3.270 -36.230 3.720 -36.160 ;
        RECT 1.420 -36.470 3.720 -36.230 ;
        RECT 1.420 -36.580 1.870 -36.470 ;
        RECT 3.270 -36.580 3.720 -36.470 ;
        RECT 4.670 -36.230 5.120 -36.130 ;
        RECT 6.520 -36.230 6.970 -36.130 ;
        RECT 4.670 -36.470 6.970 -36.230 ;
        RECT 4.670 -36.550 5.120 -36.470 ;
        RECT 5.720 -36.910 6.130 -36.470 ;
        RECT 6.520 -36.580 6.970 -36.470 ;
        RECT 8.160 -36.230 8.610 -36.130 ;
        RECT 10.010 -36.230 10.460 -36.130 ;
        RECT 8.160 -36.470 10.460 -36.230 ;
        RECT 8.160 -36.580 8.610 -36.470 ;
        RECT 9.000 -36.910 9.410 -36.470 ;
        RECT 10.010 -36.550 10.460 -36.470 ;
        RECT 11.410 -36.230 11.860 -36.160 ;
        RECT 12.460 -36.230 12.870 -35.800 ;
        RECT 13.260 -36.230 13.710 -36.130 ;
        RECT 11.410 -36.470 13.710 -36.230 ;
        RECT 11.410 -36.580 11.860 -36.470 ;
        RECT 13.260 -36.580 13.710 -36.470 ;
        RECT 14.920 -36.230 15.370 -36.130 ;
        RECT 15.760 -36.230 16.170 -35.800 ;
        RECT 18.920 -35.870 20.470 -35.650 ;
        RECT 20.850 -35.660 21.280 -35.600 ;
        RECT 21.660 -35.650 22.110 -35.600 ;
        RECT 22.710 -35.650 23.210 -35.260 ;
        RECT 21.660 -35.870 23.210 -35.650 ;
        RECT 32.420 -35.260 33.970 -35.040 ;
        RECT 32.420 -35.650 32.920 -35.260 ;
        RECT 33.520 -35.310 33.970 -35.260 ;
        RECT 34.350 -35.310 34.780 -35.250 ;
        RECT 35.160 -35.260 36.710 -35.040 ;
        RECT 39.460 -35.110 39.870 -34.680 ;
        RECT 40.260 -34.780 40.710 -34.680 ;
        RECT 41.920 -34.440 42.370 -34.330 ;
        RECT 43.770 -34.440 44.220 -34.330 ;
        RECT 41.920 -34.680 44.220 -34.440 ;
        RECT 41.920 -34.780 42.370 -34.680 ;
        RECT 42.760 -35.110 43.170 -34.680 ;
        RECT 43.770 -34.750 44.220 -34.680 ;
        RECT 45.170 -34.440 45.620 -34.360 ;
        RECT 46.220 -34.440 46.630 -34.000 ;
        RECT 47.020 -34.440 47.470 -34.330 ;
        RECT 45.170 -34.680 47.470 -34.440 ;
        RECT 45.170 -34.780 45.620 -34.680 ;
        RECT 47.020 -34.780 47.470 -34.680 ;
        RECT 48.660 -34.440 49.110 -34.330 ;
        RECT 49.500 -34.440 49.910 -34.000 ;
        RECT 52.680 -34.270 53.130 -33.990 ;
        RECT 56.500 -34.270 56.950 -33.990 ;
        RECT 66.180 -33.990 67.710 -33.780 ;
        RECT 68.090 -33.870 68.540 -33.780 ;
        RECT 68.920 -33.990 70.450 -33.780 ;
        RECT 50.510 -34.440 50.960 -34.360 ;
        RECT 48.660 -34.680 50.960 -34.440 ;
        RECT 48.660 -34.780 49.110 -34.680 ;
        RECT 50.510 -34.780 50.960 -34.680 ;
        RECT 51.910 -34.440 52.360 -34.330 ;
        RECT 53.760 -34.440 54.210 -34.330 ;
        RECT 51.910 -34.680 54.210 -34.440 ;
        RECT 51.910 -34.750 52.360 -34.680 ;
        RECT 35.160 -35.310 35.610 -35.260 ;
        RECT 33.520 -35.600 35.610 -35.310 ;
        RECT 33.520 -35.650 33.970 -35.600 ;
        RECT 16.770 -36.230 17.220 -36.160 ;
        RECT 14.920 -36.470 17.220 -36.230 ;
        RECT 14.920 -36.580 15.370 -36.470 ;
        RECT 16.770 -36.580 17.220 -36.470 ;
        RECT 18.170 -36.230 18.620 -36.130 ;
        RECT 20.020 -36.230 20.470 -36.130 ;
        RECT 18.170 -36.470 20.470 -36.230 ;
        RECT 18.170 -36.550 18.620 -36.470 ;
        RECT 12.180 -36.920 12.630 -36.640 ;
        RECT 16.000 -36.920 16.450 -36.640 ;
        RECT 19.220 -36.910 19.630 -36.470 ;
        RECT 20.020 -36.580 20.470 -36.470 ;
        RECT 21.660 -36.230 22.110 -36.130 ;
        RECT 23.510 -36.230 23.960 -36.130 ;
        RECT 21.660 -36.470 23.960 -36.230 ;
        RECT 21.660 -36.580 22.110 -36.470 ;
        RECT 22.500 -36.910 22.910 -36.470 ;
        RECT 23.510 -36.550 23.960 -36.470 ;
        RECT 24.910 -36.230 25.360 -36.160 ;
        RECT 25.960 -36.230 26.370 -35.800 ;
        RECT 26.760 -36.230 27.210 -36.130 ;
        RECT 24.910 -36.470 27.210 -36.230 ;
        RECT 24.910 -36.580 25.360 -36.470 ;
        RECT 26.760 -36.580 27.210 -36.470 ;
        RECT 28.420 -36.230 28.870 -36.130 ;
        RECT 29.260 -36.230 29.670 -35.800 ;
        RECT 32.420 -35.870 33.970 -35.650 ;
        RECT 34.350 -35.660 34.780 -35.600 ;
        RECT 35.160 -35.650 35.610 -35.600 ;
        RECT 36.210 -35.650 36.710 -35.260 ;
        RECT 35.160 -35.870 36.710 -35.650 ;
        RECT 45.920 -35.260 47.470 -35.040 ;
        RECT 45.920 -35.650 46.420 -35.260 ;
        RECT 47.020 -35.310 47.470 -35.260 ;
        RECT 47.850 -35.310 48.280 -35.250 ;
        RECT 48.660 -35.260 50.210 -35.040 ;
        RECT 52.960 -35.110 53.370 -34.680 ;
        RECT 53.760 -34.780 54.210 -34.680 ;
        RECT 55.420 -34.440 55.870 -34.330 ;
        RECT 57.270 -34.440 57.720 -34.330 ;
        RECT 55.420 -34.680 57.720 -34.440 ;
        RECT 55.420 -34.780 55.870 -34.680 ;
        RECT 56.260 -35.110 56.670 -34.680 ;
        RECT 57.270 -34.750 57.720 -34.680 ;
        RECT 58.670 -34.440 59.120 -34.360 ;
        RECT 59.720 -34.440 60.130 -34.000 ;
        RECT 60.520 -34.440 60.970 -34.330 ;
        RECT 58.670 -34.680 60.970 -34.440 ;
        RECT 58.670 -34.780 59.120 -34.680 ;
        RECT 60.520 -34.780 60.970 -34.680 ;
        RECT 62.160 -34.440 62.610 -34.330 ;
        RECT 63.000 -34.440 63.410 -34.000 ;
        RECT 66.180 -34.270 66.630 -33.990 ;
        RECT 70.000 -34.270 70.450 -33.990 ;
        RECT 79.680 -33.990 81.210 -33.780 ;
        RECT 81.590 -33.870 82.040 -33.780 ;
        RECT 82.420 -33.990 83.950 -33.780 ;
        RECT 64.010 -34.440 64.460 -34.360 ;
        RECT 62.160 -34.680 64.460 -34.440 ;
        RECT 62.160 -34.780 62.610 -34.680 ;
        RECT 64.010 -34.780 64.460 -34.680 ;
        RECT 65.410 -34.440 65.860 -34.330 ;
        RECT 67.260 -34.440 67.710 -34.330 ;
        RECT 65.410 -34.680 67.710 -34.440 ;
        RECT 65.410 -34.750 65.860 -34.680 ;
        RECT 48.660 -35.310 49.110 -35.260 ;
        RECT 47.020 -35.600 49.110 -35.310 ;
        RECT 47.020 -35.650 47.470 -35.600 ;
        RECT 30.270 -36.230 30.720 -36.160 ;
        RECT 28.420 -36.470 30.720 -36.230 ;
        RECT 28.420 -36.580 28.870 -36.470 ;
        RECT 30.270 -36.580 30.720 -36.470 ;
        RECT 31.670 -36.230 32.120 -36.130 ;
        RECT 33.520 -36.230 33.970 -36.130 ;
        RECT 31.670 -36.470 33.970 -36.230 ;
        RECT 31.670 -36.550 32.120 -36.470 ;
        RECT 12.180 -37.130 13.710 -36.920 ;
        RECT 14.090 -37.130 14.540 -37.040 ;
        RECT 14.920 -37.130 16.450 -36.920 ;
        RECT 25.680 -36.920 26.130 -36.640 ;
        RECT 29.500 -36.920 29.950 -36.640 ;
        RECT 32.720 -36.910 33.130 -36.470 ;
        RECT 33.520 -36.580 33.970 -36.470 ;
        RECT 35.160 -36.230 35.610 -36.130 ;
        RECT 37.010 -36.230 37.460 -36.130 ;
        RECT 35.160 -36.470 37.460 -36.230 ;
        RECT 35.160 -36.580 35.610 -36.470 ;
        RECT 36.000 -36.910 36.410 -36.470 ;
        RECT 37.010 -36.550 37.460 -36.470 ;
        RECT 38.410 -36.230 38.860 -36.160 ;
        RECT 39.460 -36.230 39.870 -35.800 ;
        RECT 40.260 -36.230 40.710 -36.130 ;
        RECT 38.410 -36.470 40.710 -36.230 ;
        RECT 38.410 -36.580 38.860 -36.470 ;
        RECT 40.260 -36.580 40.710 -36.470 ;
        RECT 41.920 -36.230 42.370 -36.130 ;
        RECT 42.760 -36.230 43.170 -35.800 ;
        RECT 45.920 -35.870 47.470 -35.650 ;
        RECT 47.850 -35.660 48.280 -35.600 ;
        RECT 48.660 -35.650 49.110 -35.600 ;
        RECT 49.710 -35.650 50.210 -35.260 ;
        RECT 48.660 -35.870 50.210 -35.650 ;
        RECT 59.420 -35.260 60.970 -35.040 ;
        RECT 59.420 -35.650 59.920 -35.260 ;
        RECT 60.520 -35.310 60.970 -35.260 ;
        RECT 61.350 -35.310 61.780 -35.250 ;
        RECT 62.160 -35.260 63.710 -35.040 ;
        RECT 66.460 -35.110 66.870 -34.680 ;
        RECT 67.260 -34.780 67.710 -34.680 ;
        RECT 68.920 -34.440 69.370 -34.330 ;
        RECT 70.770 -34.440 71.220 -34.330 ;
        RECT 68.920 -34.680 71.220 -34.440 ;
        RECT 68.920 -34.780 69.370 -34.680 ;
        RECT 69.760 -35.110 70.170 -34.680 ;
        RECT 70.770 -34.750 71.220 -34.680 ;
        RECT 72.170 -34.440 72.620 -34.360 ;
        RECT 73.220 -34.440 73.630 -34.000 ;
        RECT 74.020 -34.440 74.470 -34.330 ;
        RECT 72.170 -34.680 74.470 -34.440 ;
        RECT 72.170 -34.780 72.620 -34.680 ;
        RECT 74.020 -34.780 74.470 -34.680 ;
        RECT 75.660 -34.440 76.110 -34.330 ;
        RECT 76.500 -34.440 76.910 -34.000 ;
        RECT 79.680 -34.270 80.130 -33.990 ;
        RECT 83.500 -34.270 83.950 -33.990 ;
        RECT 93.180 -33.990 94.710 -33.780 ;
        RECT 95.090 -33.870 95.540 -33.780 ;
        RECT 95.920 -33.990 97.450 -33.780 ;
        RECT 77.510 -34.440 77.960 -34.360 ;
        RECT 75.660 -34.680 77.960 -34.440 ;
        RECT 75.660 -34.780 76.110 -34.680 ;
        RECT 77.510 -34.780 77.960 -34.680 ;
        RECT 78.910 -34.440 79.360 -34.330 ;
        RECT 80.760 -34.440 81.210 -34.330 ;
        RECT 78.910 -34.680 81.210 -34.440 ;
        RECT 78.910 -34.750 79.360 -34.680 ;
        RECT 62.160 -35.310 62.610 -35.260 ;
        RECT 60.520 -35.600 62.610 -35.310 ;
        RECT 60.520 -35.650 60.970 -35.600 ;
        RECT 43.770 -36.230 44.220 -36.160 ;
        RECT 41.920 -36.470 44.220 -36.230 ;
        RECT 41.920 -36.580 42.370 -36.470 ;
        RECT 43.770 -36.580 44.220 -36.470 ;
        RECT 45.170 -36.230 45.620 -36.130 ;
        RECT 47.020 -36.230 47.470 -36.130 ;
        RECT 45.170 -36.470 47.470 -36.230 ;
        RECT 45.170 -36.550 45.620 -36.470 ;
        RECT 25.680 -37.130 27.210 -36.920 ;
        RECT 27.590 -37.130 28.040 -37.040 ;
        RECT 28.420 -37.130 29.950 -36.920 ;
        RECT 39.180 -36.920 39.630 -36.640 ;
        RECT 43.000 -36.920 43.450 -36.640 ;
        RECT 46.220 -36.910 46.630 -36.470 ;
        RECT 47.020 -36.580 47.470 -36.470 ;
        RECT 48.660 -36.230 49.110 -36.130 ;
        RECT 50.510 -36.230 50.960 -36.130 ;
        RECT 48.660 -36.470 50.960 -36.230 ;
        RECT 48.660 -36.580 49.110 -36.470 ;
        RECT 49.500 -36.910 49.910 -36.470 ;
        RECT 50.510 -36.550 50.960 -36.470 ;
        RECT 51.910 -36.230 52.360 -36.160 ;
        RECT 52.960 -36.230 53.370 -35.800 ;
        RECT 53.760 -36.230 54.210 -36.130 ;
        RECT 51.910 -36.470 54.210 -36.230 ;
        RECT 51.910 -36.580 52.360 -36.470 ;
        RECT 53.760 -36.580 54.210 -36.470 ;
        RECT 55.420 -36.230 55.870 -36.130 ;
        RECT 56.260 -36.230 56.670 -35.800 ;
        RECT 59.420 -35.870 60.970 -35.650 ;
        RECT 61.350 -35.660 61.780 -35.600 ;
        RECT 62.160 -35.650 62.610 -35.600 ;
        RECT 63.210 -35.650 63.710 -35.260 ;
        RECT 62.160 -35.870 63.710 -35.650 ;
        RECT 72.920 -35.260 74.470 -35.040 ;
        RECT 72.920 -35.650 73.420 -35.260 ;
        RECT 74.020 -35.310 74.470 -35.260 ;
        RECT 74.850 -35.310 75.280 -35.250 ;
        RECT 75.660 -35.260 77.210 -35.040 ;
        RECT 79.960 -35.110 80.370 -34.680 ;
        RECT 80.760 -34.780 81.210 -34.680 ;
        RECT 82.420 -34.440 82.870 -34.330 ;
        RECT 84.270 -34.440 84.720 -34.330 ;
        RECT 82.420 -34.680 84.720 -34.440 ;
        RECT 82.420 -34.780 82.870 -34.680 ;
        RECT 83.260 -35.110 83.670 -34.680 ;
        RECT 84.270 -34.750 84.720 -34.680 ;
        RECT 85.670 -34.440 86.120 -34.360 ;
        RECT 86.720 -34.440 87.130 -34.000 ;
        RECT 87.520 -34.440 87.970 -34.330 ;
        RECT 85.670 -34.680 87.970 -34.440 ;
        RECT 85.670 -34.780 86.120 -34.680 ;
        RECT 87.520 -34.780 87.970 -34.680 ;
        RECT 89.160 -34.440 89.610 -34.330 ;
        RECT 90.000 -34.440 90.410 -34.000 ;
        RECT 93.180 -34.270 93.630 -33.990 ;
        RECT 97.000 -34.270 97.450 -33.990 ;
        RECT 106.680 -33.990 108.210 -33.780 ;
        RECT 108.590 -33.870 109.040 -33.780 ;
        RECT 109.420 -33.990 110.950 -33.780 ;
        RECT 91.010 -34.440 91.460 -34.360 ;
        RECT 89.160 -34.680 91.460 -34.440 ;
        RECT 89.160 -34.780 89.610 -34.680 ;
        RECT 91.010 -34.780 91.460 -34.680 ;
        RECT 92.410 -34.440 92.860 -34.330 ;
        RECT 94.260 -34.440 94.710 -34.330 ;
        RECT 92.410 -34.680 94.710 -34.440 ;
        RECT 92.410 -34.750 92.860 -34.680 ;
        RECT 75.660 -35.310 76.110 -35.260 ;
        RECT 74.020 -35.600 76.110 -35.310 ;
        RECT 74.020 -35.650 74.470 -35.600 ;
        RECT 57.270 -36.230 57.720 -36.160 ;
        RECT 55.420 -36.470 57.720 -36.230 ;
        RECT 55.420 -36.580 55.870 -36.470 ;
        RECT 57.270 -36.580 57.720 -36.470 ;
        RECT 58.670 -36.230 59.120 -36.130 ;
        RECT 60.520 -36.230 60.970 -36.130 ;
        RECT 58.670 -36.470 60.970 -36.230 ;
        RECT 58.670 -36.550 59.120 -36.470 ;
        RECT 39.180 -37.130 40.710 -36.920 ;
        RECT 41.090 -37.130 41.540 -37.040 ;
        RECT 41.920 -37.130 43.450 -36.920 ;
        RECT 52.680 -36.920 53.130 -36.640 ;
        RECT 56.500 -36.920 56.950 -36.640 ;
        RECT 59.720 -36.910 60.130 -36.470 ;
        RECT 60.520 -36.580 60.970 -36.470 ;
        RECT 62.160 -36.230 62.610 -36.130 ;
        RECT 64.010 -36.230 64.460 -36.130 ;
        RECT 62.160 -36.470 64.460 -36.230 ;
        RECT 62.160 -36.580 62.610 -36.470 ;
        RECT 63.000 -36.910 63.410 -36.470 ;
        RECT 64.010 -36.550 64.460 -36.470 ;
        RECT 65.410 -36.230 65.860 -36.160 ;
        RECT 66.460 -36.230 66.870 -35.800 ;
        RECT 67.260 -36.230 67.710 -36.130 ;
        RECT 65.410 -36.470 67.710 -36.230 ;
        RECT 65.410 -36.580 65.860 -36.470 ;
        RECT 67.260 -36.580 67.710 -36.470 ;
        RECT 68.920 -36.230 69.370 -36.130 ;
        RECT 69.760 -36.230 70.170 -35.800 ;
        RECT 72.920 -35.870 74.470 -35.650 ;
        RECT 74.850 -35.660 75.280 -35.600 ;
        RECT 75.660 -35.650 76.110 -35.600 ;
        RECT 76.710 -35.650 77.210 -35.260 ;
        RECT 75.660 -35.870 77.210 -35.650 ;
        RECT 86.420 -35.260 87.970 -35.040 ;
        RECT 86.420 -35.650 86.920 -35.260 ;
        RECT 87.520 -35.310 87.970 -35.260 ;
        RECT 88.350 -35.310 88.780 -35.250 ;
        RECT 89.160 -35.260 90.710 -35.040 ;
        RECT 93.460 -35.110 93.870 -34.680 ;
        RECT 94.260 -34.780 94.710 -34.680 ;
        RECT 95.920 -34.440 96.370 -34.330 ;
        RECT 97.770 -34.440 98.220 -34.330 ;
        RECT 95.920 -34.680 98.220 -34.440 ;
        RECT 95.920 -34.780 96.370 -34.680 ;
        RECT 96.760 -35.110 97.170 -34.680 ;
        RECT 97.770 -34.750 98.220 -34.680 ;
        RECT 99.170 -34.440 99.620 -34.360 ;
        RECT 100.220 -34.440 100.630 -34.000 ;
        RECT 101.020 -34.440 101.470 -34.330 ;
        RECT 99.170 -34.680 101.470 -34.440 ;
        RECT 99.170 -34.780 99.620 -34.680 ;
        RECT 101.020 -34.780 101.470 -34.680 ;
        RECT 102.660 -34.440 103.110 -34.330 ;
        RECT 103.500 -34.440 103.910 -34.000 ;
        RECT 106.680 -34.270 107.130 -33.990 ;
        RECT 110.500 -34.270 110.950 -33.990 ;
        RECT 120.180 -33.990 121.710 -33.780 ;
        RECT 122.090 -33.870 122.540 -33.780 ;
        RECT 122.920 -33.990 124.450 -33.780 ;
        RECT 104.510 -34.440 104.960 -34.360 ;
        RECT 102.660 -34.680 104.960 -34.440 ;
        RECT 102.660 -34.780 103.110 -34.680 ;
        RECT 104.510 -34.780 104.960 -34.680 ;
        RECT 105.910 -34.440 106.360 -34.330 ;
        RECT 107.760 -34.440 108.210 -34.330 ;
        RECT 105.910 -34.680 108.210 -34.440 ;
        RECT 105.910 -34.750 106.360 -34.680 ;
        RECT 89.160 -35.310 89.610 -35.260 ;
        RECT 87.520 -35.600 89.610 -35.310 ;
        RECT 87.520 -35.650 87.970 -35.600 ;
        RECT 70.770 -36.230 71.220 -36.160 ;
        RECT 68.920 -36.470 71.220 -36.230 ;
        RECT 68.920 -36.580 69.370 -36.470 ;
        RECT 70.770 -36.580 71.220 -36.470 ;
        RECT 72.170 -36.230 72.620 -36.130 ;
        RECT 74.020 -36.230 74.470 -36.130 ;
        RECT 72.170 -36.470 74.470 -36.230 ;
        RECT 72.170 -36.550 72.620 -36.470 ;
        RECT 52.680 -37.130 54.210 -36.920 ;
        RECT 54.590 -37.130 55.040 -37.040 ;
        RECT 55.420 -37.130 56.950 -36.920 ;
        RECT 66.180 -36.920 66.630 -36.640 ;
        RECT 70.000 -36.920 70.450 -36.640 ;
        RECT 73.220 -36.910 73.630 -36.470 ;
        RECT 74.020 -36.580 74.470 -36.470 ;
        RECT 75.660 -36.230 76.110 -36.130 ;
        RECT 77.510 -36.230 77.960 -36.130 ;
        RECT 75.660 -36.470 77.960 -36.230 ;
        RECT 75.660 -36.580 76.110 -36.470 ;
        RECT 76.500 -36.910 76.910 -36.470 ;
        RECT 77.510 -36.550 77.960 -36.470 ;
        RECT 78.910 -36.230 79.360 -36.160 ;
        RECT 79.960 -36.230 80.370 -35.800 ;
        RECT 80.760 -36.230 81.210 -36.130 ;
        RECT 78.910 -36.470 81.210 -36.230 ;
        RECT 78.910 -36.580 79.360 -36.470 ;
        RECT 80.760 -36.580 81.210 -36.470 ;
        RECT 82.420 -36.230 82.870 -36.130 ;
        RECT 83.260 -36.230 83.670 -35.800 ;
        RECT 86.420 -35.870 87.970 -35.650 ;
        RECT 88.350 -35.660 88.780 -35.600 ;
        RECT 89.160 -35.650 89.610 -35.600 ;
        RECT 90.210 -35.650 90.710 -35.260 ;
        RECT 89.160 -35.870 90.710 -35.650 ;
        RECT 99.920 -35.260 101.470 -35.040 ;
        RECT 99.920 -35.650 100.420 -35.260 ;
        RECT 101.020 -35.310 101.470 -35.260 ;
        RECT 101.850 -35.310 102.280 -35.250 ;
        RECT 102.660 -35.260 104.210 -35.040 ;
        RECT 106.960 -35.110 107.370 -34.680 ;
        RECT 107.760 -34.780 108.210 -34.680 ;
        RECT 109.420 -34.440 109.870 -34.330 ;
        RECT 111.270 -34.440 111.720 -34.330 ;
        RECT 109.420 -34.680 111.720 -34.440 ;
        RECT 109.420 -34.780 109.870 -34.680 ;
        RECT 110.260 -35.110 110.670 -34.680 ;
        RECT 111.270 -34.750 111.720 -34.680 ;
        RECT 112.670 -34.440 113.120 -34.360 ;
        RECT 113.720 -34.440 114.130 -34.000 ;
        RECT 114.520 -34.440 114.970 -34.330 ;
        RECT 112.670 -34.680 114.970 -34.440 ;
        RECT 112.670 -34.780 113.120 -34.680 ;
        RECT 114.520 -34.780 114.970 -34.680 ;
        RECT 116.160 -34.440 116.610 -34.330 ;
        RECT 117.000 -34.440 117.410 -34.000 ;
        RECT 120.180 -34.270 120.630 -33.990 ;
        RECT 124.000 -34.270 124.450 -33.990 ;
        RECT 133.680 -33.990 135.210 -33.780 ;
        RECT 135.590 -33.870 136.040 -33.780 ;
        RECT 136.420 -33.990 137.950 -33.780 ;
        RECT 118.010 -34.440 118.460 -34.360 ;
        RECT 116.160 -34.680 118.460 -34.440 ;
        RECT 116.160 -34.780 116.610 -34.680 ;
        RECT 118.010 -34.780 118.460 -34.680 ;
        RECT 119.410 -34.440 119.860 -34.330 ;
        RECT 121.260 -34.440 121.710 -34.330 ;
        RECT 119.410 -34.680 121.710 -34.440 ;
        RECT 119.410 -34.750 119.860 -34.680 ;
        RECT 102.660 -35.310 103.110 -35.260 ;
        RECT 101.020 -35.600 103.110 -35.310 ;
        RECT 101.020 -35.650 101.470 -35.600 ;
        RECT 84.270 -36.230 84.720 -36.160 ;
        RECT 82.420 -36.470 84.720 -36.230 ;
        RECT 82.420 -36.580 82.870 -36.470 ;
        RECT 84.270 -36.580 84.720 -36.470 ;
        RECT 85.670 -36.230 86.120 -36.130 ;
        RECT 87.520 -36.230 87.970 -36.130 ;
        RECT 85.670 -36.470 87.970 -36.230 ;
        RECT 85.670 -36.550 86.120 -36.470 ;
        RECT 66.180 -37.130 67.710 -36.920 ;
        RECT 68.090 -37.130 68.540 -37.040 ;
        RECT 68.920 -37.130 70.450 -36.920 ;
        RECT 79.680 -36.920 80.130 -36.640 ;
        RECT 83.500 -36.920 83.950 -36.640 ;
        RECT 86.720 -36.910 87.130 -36.470 ;
        RECT 87.520 -36.580 87.970 -36.470 ;
        RECT 89.160 -36.230 89.610 -36.130 ;
        RECT 91.010 -36.230 91.460 -36.130 ;
        RECT 89.160 -36.470 91.460 -36.230 ;
        RECT 89.160 -36.580 89.610 -36.470 ;
        RECT 90.000 -36.910 90.410 -36.470 ;
        RECT 91.010 -36.550 91.460 -36.470 ;
        RECT 92.410 -36.230 92.860 -36.160 ;
        RECT 93.460 -36.230 93.870 -35.800 ;
        RECT 94.260 -36.230 94.710 -36.130 ;
        RECT 92.410 -36.470 94.710 -36.230 ;
        RECT 92.410 -36.580 92.860 -36.470 ;
        RECT 94.260 -36.580 94.710 -36.470 ;
        RECT 95.920 -36.230 96.370 -36.130 ;
        RECT 96.760 -36.230 97.170 -35.800 ;
        RECT 99.920 -35.870 101.470 -35.650 ;
        RECT 101.850 -35.660 102.280 -35.600 ;
        RECT 102.660 -35.650 103.110 -35.600 ;
        RECT 103.710 -35.650 104.210 -35.260 ;
        RECT 102.660 -35.870 104.210 -35.650 ;
        RECT 113.420 -35.260 114.970 -35.040 ;
        RECT 113.420 -35.650 113.920 -35.260 ;
        RECT 114.520 -35.310 114.970 -35.260 ;
        RECT 115.350 -35.310 115.780 -35.250 ;
        RECT 116.160 -35.260 117.710 -35.040 ;
        RECT 120.460 -35.110 120.870 -34.680 ;
        RECT 121.260 -34.780 121.710 -34.680 ;
        RECT 122.920 -34.440 123.370 -34.330 ;
        RECT 124.770 -34.440 125.220 -34.330 ;
        RECT 122.920 -34.680 125.220 -34.440 ;
        RECT 122.920 -34.780 123.370 -34.680 ;
        RECT 123.760 -35.110 124.170 -34.680 ;
        RECT 124.770 -34.750 125.220 -34.680 ;
        RECT 126.170 -34.440 126.620 -34.360 ;
        RECT 127.220 -34.440 127.630 -34.000 ;
        RECT 128.020 -34.440 128.470 -34.330 ;
        RECT 126.170 -34.680 128.470 -34.440 ;
        RECT 126.170 -34.780 126.620 -34.680 ;
        RECT 128.020 -34.780 128.470 -34.680 ;
        RECT 129.660 -34.440 130.110 -34.330 ;
        RECT 130.500 -34.440 130.910 -34.000 ;
        RECT 133.680 -34.270 134.130 -33.990 ;
        RECT 137.500 -34.270 137.950 -33.990 ;
        RECT 147.180 -33.990 148.710 -33.780 ;
        RECT 149.090 -33.870 149.540 -33.780 ;
        RECT 149.920 -33.990 151.450 -33.780 ;
        RECT 131.510 -34.440 131.960 -34.360 ;
        RECT 129.660 -34.680 131.960 -34.440 ;
        RECT 129.660 -34.780 130.110 -34.680 ;
        RECT 131.510 -34.780 131.960 -34.680 ;
        RECT 132.910 -34.440 133.360 -34.330 ;
        RECT 134.760 -34.440 135.210 -34.330 ;
        RECT 132.910 -34.680 135.210 -34.440 ;
        RECT 132.910 -34.750 133.360 -34.680 ;
        RECT 116.160 -35.310 116.610 -35.260 ;
        RECT 114.520 -35.600 116.610 -35.310 ;
        RECT 114.520 -35.650 114.970 -35.600 ;
        RECT 97.770 -36.230 98.220 -36.160 ;
        RECT 95.920 -36.470 98.220 -36.230 ;
        RECT 95.920 -36.580 96.370 -36.470 ;
        RECT 97.770 -36.580 98.220 -36.470 ;
        RECT 99.170 -36.230 99.620 -36.130 ;
        RECT 101.020 -36.230 101.470 -36.130 ;
        RECT 99.170 -36.470 101.470 -36.230 ;
        RECT 99.170 -36.550 99.620 -36.470 ;
        RECT 79.680 -37.130 81.210 -36.920 ;
        RECT 81.590 -37.130 82.040 -37.040 ;
        RECT 82.420 -37.130 83.950 -36.920 ;
        RECT 93.180 -36.920 93.630 -36.640 ;
        RECT 97.000 -36.920 97.450 -36.640 ;
        RECT 100.220 -36.910 100.630 -36.470 ;
        RECT 101.020 -36.580 101.470 -36.470 ;
        RECT 102.660 -36.230 103.110 -36.130 ;
        RECT 104.510 -36.230 104.960 -36.130 ;
        RECT 102.660 -36.470 104.960 -36.230 ;
        RECT 102.660 -36.580 103.110 -36.470 ;
        RECT 103.500 -36.910 103.910 -36.470 ;
        RECT 104.510 -36.550 104.960 -36.470 ;
        RECT 105.910 -36.230 106.360 -36.160 ;
        RECT 106.960 -36.230 107.370 -35.800 ;
        RECT 107.760 -36.230 108.210 -36.130 ;
        RECT 105.910 -36.470 108.210 -36.230 ;
        RECT 105.910 -36.580 106.360 -36.470 ;
        RECT 107.760 -36.580 108.210 -36.470 ;
        RECT 109.420 -36.230 109.870 -36.130 ;
        RECT 110.260 -36.230 110.670 -35.800 ;
        RECT 113.420 -35.870 114.970 -35.650 ;
        RECT 115.350 -35.660 115.780 -35.600 ;
        RECT 116.160 -35.650 116.610 -35.600 ;
        RECT 117.210 -35.650 117.710 -35.260 ;
        RECT 116.160 -35.870 117.710 -35.650 ;
        RECT 126.920 -35.260 128.470 -35.040 ;
        RECT 126.920 -35.650 127.420 -35.260 ;
        RECT 128.020 -35.310 128.470 -35.260 ;
        RECT 128.850 -35.310 129.280 -35.250 ;
        RECT 129.660 -35.260 131.210 -35.040 ;
        RECT 133.960 -35.110 134.370 -34.680 ;
        RECT 134.760 -34.780 135.210 -34.680 ;
        RECT 136.420 -34.440 136.870 -34.330 ;
        RECT 138.270 -34.440 138.720 -34.330 ;
        RECT 136.420 -34.680 138.720 -34.440 ;
        RECT 136.420 -34.780 136.870 -34.680 ;
        RECT 137.260 -35.110 137.670 -34.680 ;
        RECT 138.270 -34.750 138.720 -34.680 ;
        RECT 139.670 -34.440 140.120 -34.360 ;
        RECT 140.720 -34.440 141.130 -34.000 ;
        RECT 141.520 -34.440 141.970 -34.330 ;
        RECT 139.670 -34.680 141.970 -34.440 ;
        RECT 139.670 -34.780 140.120 -34.680 ;
        RECT 141.520 -34.780 141.970 -34.680 ;
        RECT 143.160 -34.440 143.610 -34.330 ;
        RECT 144.000 -34.440 144.410 -34.000 ;
        RECT 147.180 -34.270 147.630 -33.990 ;
        RECT 151.000 -34.270 151.450 -33.990 ;
        RECT 160.680 -33.990 162.210 -33.780 ;
        RECT 162.590 -33.870 163.040 -33.780 ;
        RECT 163.420 -33.990 164.950 -33.780 ;
        RECT 145.010 -34.440 145.460 -34.360 ;
        RECT 143.160 -34.680 145.460 -34.440 ;
        RECT 143.160 -34.780 143.610 -34.680 ;
        RECT 145.010 -34.780 145.460 -34.680 ;
        RECT 146.410 -34.440 146.860 -34.330 ;
        RECT 148.260 -34.440 148.710 -34.330 ;
        RECT 146.410 -34.680 148.710 -34.440 ;
        RECT 146.410 -34.750 146.860 -34.680 ;
        RECT 129.660 -35.310 130.110 -35.260 ;
        RECT 128.020 -35.600 130.110 -35.310 ;
        RECT 128.020 -35.650 128.470 -35.600 ;
        RECT 111.270 -36.230 111.720 -36.160 ;
        RECT 109.420 -36.470 111.720 -36.230 ;
        RECT 109.420 -36.580 109.870 -36.470 ;
        RECT 111.270 -36.580 111.720 -36.470 ;
        RECT 112.670 -36.230 113.120 -36.130 ;
        RECT 114.520 -36.230 114.970 -36.130 ;
        RECT 112.670 -36.470 114.970 -36.230 ;
        RECT 112.670 -36.550 113.120 -36.470 ;
        RECT 93.180 -37.130 94.710 -36.920 ;
        RECT 95.090 -37.130 95.540 -37.040 ;
        RECT 95.920 -37.130 97.450 -36.920 ;
        RECT 106.680 -36.920 107.130 -36.640 ;
        RECT 110.500 -36.920 110.950 -36.640 ;
        RECT 113.720 -36.910 114.130 -36.470 ;
        RECT 114.520 -36.580 114.970 -36.470 ;
        RECT 116.160 -36.230 116.610 -36.130 ;
        RECT 118.010 -36.230 118.460 -36.130 ;
        RECT 116.160 -36.470 118.460 -36.230 ;
        RECT 116.160 -36.580 116.610 -36.470 ;
        RECT 117.000 -36.910 117.410 -36.470 ;
        RECT 118.010 -36.550 118.460 -36.470 ;
        RECT 119.410 -36.230 119.860 -36.160 ;
        RECT 120.460 -36.230 120.870 -35.800 ;
        RECT 121.260 -36.230 121.710 -36.130 ;
        RECT 119.410 -36.470 121.710 -36.230 ;
        RECT 119.410 -36.580 119.860 -36.470 ;
        RECT 121.260 -36.580 121.710 -36.470 ;
        RECT 122.920 -36.230 123.370 -36.130 ;
        RECT 123.760 -36.230 124.170 -35.800 ;
        RECT 126.920 -35.870 128.470 -35.650 ;
        RECT 128.850 -35.660 129.280 -35.600 ;
        RECT 129.660 -35.650 130.110 -35.600 ;
        RECT 130.710 -35.650 131.210 -35.260 ;
        RECT 129.660 -35.870 131.210 -35.650 ;
        RECT 140.420 -35.260 141.970 -35.040 ;
        RECT 140.420 -35.650 140.920 -35.260 ;
        RECT 141.520 -35.310 141.970 -35.260 ;
        RECT 142.350 -35.310 142.780 -35.250 ;
        RECT 143.160 -35.260 144.710 -35.040 ;
        RECT 147.460 -35.110 147.870 -34.680 ;
        RECT 148.260 -34.780 148.710 -34.680 ;
        RECT 149.920 -34.440 150.370 -34.330 ;
        RECT 151.770 -34.440 152.220 -34.330 ;
        RECT 149.920 -34.680 152.220 -34.440 ;
        RECT 149.920 -34.780 150.370 -34.680 ;
        RECT 150.760 -35.110 151.170 -34.680 ;
        RECT 151.770 -34.750 152.220 -34.680 ;
        RECT 153.170 -34.440 153.620 -34.360 ;
        RECT 154.220 -34.440 154.630 -34.000 ;
        RECT 155.020 -34.440 155.470 -34.330 ;
        RECT 153.170 -34.680 155.470 -34.440 ;
        RECT 153.170 -34.780 153.620 -34.680 ;
        RECT 155.020 -34.780 155.470 -34.680 ;
        RECT 156.660 -34.440 157.110 -34.330 ;
        RECT 157.500 -34.440 157.910 -34.000 ;
        RECT 160.680 -34.270 161.130 -33.990 ;
        RECT 164.500 -34.270 164.950 -33.990 ;
        RECT 174.180 -33.990 175.710 -33.780 ;
        RECT 176.090 -33.870 176.540 -33.780 ;
        RECT 176.920 -33.990 178.450 -33.780 ;
        RECT 158.510 -34.440 158.960 -34.360 ;
        RECT 156.660 -34.680 158.960 -34.440 ;
        RECT 156.660 -34.780 157.110 -34.680 ;
        RECT 158.510 -34.780 158.960 -34.680 ;
        RECT 159.910 -34.440 160.360 -34.330 ;
        RECT 161.760 -34.440 162.210 -34.330 ;
        RECT 159.910 -34.680 162.210 -34.440 ;
        RECT 159.910 -34.750 160.360 -34.680 ;
        RECT 143.160 -35.310 143.610 -35.260 ;
        RECT 141.520 -35.600 143.610 -35.310 ;
        RECT 141.520 -35.650 141.970 -35.600 ;
        RECT 124.770 -36.230 125.220 -36.160 ;
        RECT 122.920 -36.470 125.220 -36.230 ;
        RECT 122.920 -36.580 123.370 -36.470 ;
        RECT 124.770 -36.580 125.220 -36.470 ;
        RECT 126.170 -36.230 126.620 -36.130 ;
        RECT 128.020 -36.230 128.470 -36.130 ;
        RECT 126.170 -36.470 128.470 -36.230 ;
        RECT 126.170 -36.550 126.620 -36.470 ;
        RECT 106.680 -37.130 108.210 -36.920 ;
        RECT 108.590 -37.130 109.040 -37.040 ;
        RECT 109.420 -37.130 110.950 -36.920 ;
        RECT 120.180 -36.920 120.630 -36.640 ;
        RECT 124.000 -36.920 124.450 -36.640 ;
        RECT 127.220 -36.910 127.630 -36.470 ;
        RECT 128.020 -36.580 128.470 -36.470 ;
        RECT 129.660 -36.230 130.110 -36.130 ;
        RECT 131.510 -36.230 131.960 -36.130 ;
        RECT 129.660 -36.470 131.960 -36.230 ;
        RECT 129.660 -36.580 130.110 -36.470 ;
        RECT 130.500 -36.910 130.910 -36.470 ;
        RECT 131.510 -36.550 131.960 -36.470 ;
        RECT 132.910 -36.230 133.360 -36.160 ;
        RECT 133.960 -36.230 134.370 -35.800 ;
        RECT 134.760 -36.230 135.210 -36.130 ;
        RECT 132.910 -36.470 135.210 -36.230 ;
        RECT 132.910 -36.580 133.360 -36.470 ;
        RECT 134.760 -36.580 135.210 -36.470 ;
        RECT 136.420 -36.230 136.870 -36.130 ;
        RECT 137.260 -36.230 137.670 -35.800 ;
        RECT 140.420 -35.870 141.970 -35.650 ;
        RECT 142.350 -35.660 142.780 -35.600 ;
        RECT 143.160 -35.650 143.610 -35.600 ;
        RECT 144.210 -35.650 144.710 -35.260 ;
        RECT 143.160 -35.870 144.710 -35.650 ;
        RECT 153.920 -35.260 155.470 -35.040 ;
        RECT 153.920 -35.650 154.420 -35.260 ;
        RECT 155.020 -35.310 155.470 -35.260 ;
        RECT 155.850 -35.310 156.280 -35.250 ;
        RECT 156.660 -35.260 158.210 -35.040 ;
        RECT 160.960 -35.110 161.370 -34.680 ;
        RECT 161.760 -34.780 162.210 -34.680 ;
        RECT 163.420 -34.440 163.870 -34.330 ;
        RECT 165.270 -34.440 165.720 -34.330 ;
        RECT 163.420 -34.680 165.720 -34.440 ;
        RECT 163.420 -34.780 163.870 -34.680 ;
        RECT 164.260 -35.110 164.670 -34.680 ;
        RECT 165.270 -34.750 165.720 -34.680 ;
        RECT 166.670 -34.440 167.120 -34.360 ;
        RECT 167.720 -34.440 168.130 -34.000 ;
        RECT 168.520 -34.440 168.970 -34.330 ;
        RECT 166.670 -34.680 168.970 -34.440 ;
        RECT 166.670 -34.780 167.120 -34.680 ;
        RECT 168.520 -34.780 168.970 -34.680 ;
        RECT 170.160 -34.440 170.610 -34.330 ;
        RECT 171.000 -34.440 171.410 -34.000 ;
        RECT 174.180 -34.270 174.630 -33.990 ;
        RECT 178.000 -34.270 178.450 -33.990 ;
        RECT 187.680 -33.990 189.210 -33.780 ;
        RECT 189.590 -33.870 190.040 -33.780 ;
        RECT 190.420 -33.990 191.950 -33.780 ;
        RECT 172.010 -34.440 172.460 -34.360 ;
        RECT 170.160 -34.680 172.460 -34.440 ;
        RECT 170.160 -34.780 170.610 -34.680 ;
        RECT 172.010 -34.780 172.460 -34.680 ;
        RECT 173.410 -34.440 173.860 -34.330 ;
        RECT 175.260 -34.440 175.710 -34.330 ;
        RECT 173.410 -34.680 175.710 -34.440 ;
        RECT 173.410 -34.750 173.860 -34.680 ;
        RECT 156.660 -35.310 157.110 -35.260 ;
        RECT 155.020 -35.600 157.110 -35.310 ;
        RECT 155.020 -35.650 155.470 -35.600 ;
        RECT 138.270 -36.230 138.720 -36.160 ;
        RECT 136.420 -36.470 138.720 -36.230 ;
        RECT 136.420 -36.580 136.870 -36.470 ;
        RECT 138.270 -36.580 138.720 -36.470 ;
        RECT 139.670 -36.230 140.120 -36.130 ;
        RECT 141.520 -36.230 141.970 -36.130 ;
        RECT 139.670 -36.470 141.970 -36.230 ;
        RECT 139.670 -36.550 140.120 -36.470 ;
        RECT 120.180 -37.130 121.710 -36.920 ;
        RECT 122.090 -37.130 122.540 -37.040 ;
        RECT 122.920 -37.130 124.450 -36.920 ;
        RECT 133.680 -36.920 134.130 -36.640 ;
        RECT 137.500 -36.920 137.950 -36.640 ;
        RECT 140.720 -36.910 141.130 -36.470 ;
        RECT 141.520 -36.580 141.970 -36.470 ;
        RECT 143.160 -36.230 143.610 -36.130 ;
        RECT 145.010 -36.230 145.460 -36.130 ;
        RECT 143.160 -36.470 145.460 -36.230 ;
        RECT 143.160 -36.580 143.610 -36.470 ;
        RECT 144.000 -36.910 144.410 -36.470 ;
        RECT 145.010 -36.550 145.460 -36.470 ;
        RECT 146.410 -36.230 146.860 -36.160 ;
        RECT 147.460 -36.230 147.870 -35.800 ;
        RECT 148.260 -36.230 148.710 -36.130 ;
        RECT 146.410 -36.470 148.710 -36.230 ;
        RECT 146.410 -36.580 146.860 -36.470 ;
        RECT 148.260 -36.580 148.710 -36.470 ;
        RECT 149.920 -36.230 150.370 -36.130 ;
        RECT 150.760 -36.230 151.170 -35.800 ;
        RECT 153.920 -35.870 155.470 -35.650 ;
        RECT 155.850 -35.660 156.280 -35.600 ;
        RECT 156.660 -35.650 157.110 -35.600 ;
        RECT 157.710 -35.650 158.210 -35.260 ;
        RECT 156.660 -35.870 158.210 -35.650 ;
        RECT 167.420 -35.260 168.970 -35.040 ;
        RECT 167.420 -35.650 167.920 -35.260 ;
        RECT 168.520 -35.310 168.970 -35.260 ;
        RECT 169.350 -35.310 169.780 -35.250 ;
        RECT 170.160 -35.260 171.710 -35.040 ;
        RECT 174.460 -35.110 174.870 -34.680 ;
        RECT 175.260 -34.780 175.710 -34.680 ;
        RECT 176.920 -34.440 177.370 -34.330 ;
        RECT 178.770 -34.440 179.220 -34.330 ;
        RECT 176.920 -34.680 179.220 -34.440 ;
        RECT 176.920 -34.780 177.370 -34.680 ;
        RECT 177.760 -35.110 178.170 -34.680 ;
        RECT 178.770 -34.750 179.220 -34.680 ;
        RECT 180.170 -34.440 180.620 -34.360 ;
        RECT 181.220 -34.440 181.630 -34.000 ;
        RECT 182.020 -34.440 182.470 -34.330 ;
        RECT 180.170 -34.680 182.470 -34.440 ;
        RECT 180.170 -34.780 180.620 -34.680 ;
        RECT 182.020 -34.780 182.470 -34.680 ;
        RECT 183.660 -34.440 184.110 -34.330 ;
        RECT 184.500 -34.440 184.910 -34.000 ;
        RECT 187.680 -34.270 188.130 -33.990 ;
        RECT 191.500 -34.270 191.950 -33.990 ;
        RECT 201.180 -33.990 202.710 -33.780 ;
        RECT 203.090 -33.870 203.540 -33.780 ;
        RECT 203.920 -33.990 205.450 -33.780 ;
        RECT 185.510 -34.440 185.960 -34.360 ;
        RECT 183.660 -34.680 185.960 -34.440 ;
        RECT 183.660 -34.780 184.110 -34.680 ;
        RECT 185.510 -34.780 185.960 -34.680 ;
        RECT 186.910 -34.440 187.360 -34.330 ;
        RECT 188.760 -34.440 189.210 -34.330 ;
        RECT 186.910 -34.680 189.210 -34.440 ;
        RECT 186.910 -34.750 187.360 -34.680 ;
        RECT 170.160 -35.310 170.610 -35.260 ;
        RECT 168.520 -35.600 170.610 -35.310 ;
        RECT 168.520 -35.650 168.970 -35.600 ;
        RECT 151.770 -36.230 152.220 -36.160 ;
        RECT 149.920 -36.470 152.220 -36.230 ;
        RECT 149.920 -36.580 150.370 -36.470 ;
        RECT 151.770 -36.580 152.220 -36.470 ;
        RECT 153.170 -36.230 153.620 -36.130 ;
        RECT 155.020 -36.230 155.470 -36.130 ;
        RECT 153.170 -36.470 155.470 -36.230 ;
        RECT 153.170 -36.550 153.620 -36.470 ;
        RECT 133.680 -37.130 135.210 -36.920 ;
        RECT 135.590 -37.130 136.040 -37.040 ;
        RECT 136.420 -37.130 137.950 -36.920 ;
        RECT 147.180 -36.920 147.630 -36.640 ;
        RECT 151.000 -36.920 151.450 -36.640 ;
        RECT 154.220 -36.910 154.630 -36.470 ;
        RECT 155.020 -36.580 155.470 -36.470 ;
        RECT 156.660 -36.230 157.110 -36.130 ;
        RECT 158.510 -36.230 158.960 -36.130 ;
        RECT 156.660 -36.470 158.960 -36.230 ;
        RECT 156.660 -36.580 157.110 -36.470 ;
        RECT 157.500 -36.910 157.910 -36.470 ;
        RECT 158.510 -36.550 158.960 -36.470 ;
        RECT 159.910 -36.230 160.360 -36.160 ;
        RECT 160.960 -36.230 161.370 -35.800 ;
        RECT 161.760 -36.230 162.210 -36.130 ;
        RECT 159.910 -36.470 162.210 -36.230 ;
        RECT 159.910 -36.580 160.360 -36.470 ;
        RECT 161.760 -36.580 162.210 -36.470 ;
        RECT 163.420 -36.230 163.870 -36.130 ;
        RECT 164.260 -36.230 164.670 -35.800 ;
        RECT 167.420 -35.870 168.970 -35.650 ;
        RECT 169.350 -35.660 169.780 -35.600 ;
        RECT 170.160 -35.650 170.610 -35.600 ;
        RECT 171.210 -35.650 171.710 -35.260 ;
        RECT 170.160 -35.870 171.710 -35.650 ;
        RECT 180.920 -35.260 182.470 -35.040 ;
        RECT 180.920 -35.650 181.420 -35.260 ;
        RECT 182.020 -35.310 182.470 -35.260 ;
        RECT 182.850 -35.310 183.280 -35.250 ;
        RECT 183.660 -35.260 185.210 -35.040 ;
        RECT 187.960 -35.110 188.370 -34.680 ;
        RECT 188.760 -34.780 189.210 -34.680 ;
        RECT 190.420 -34.440 190.870 -34.330 ;
        RECT 192.270 -34.440 192.720 -34.330 ;
        RECT 190.420 -34.680 192.720 -34.440 ;
        RECT 190.420 -34.780 190.870 -34.680 ;
        RECT 191.260 -35.110 191.670 -34.680 ;
        RECT 192.270 -34.750 192.720 -34.680 ;
        RECT 193.670 -34.440 194.120 -34.360 ;
        RECT 194.720 -34.440 195.130 -34.000 ;
        RECT 195.520 -34.440 195.970 -34.330 ;
        RECT 193.670 -34.680 195.970 -34.440 ;
        RECT 193.670 -34.780 194.120 -34.680 ;
        RECT 195.520 -34.780 195.970 -34.680 ;
        RECT 197.160 -34.440 197.610 -34.330 ;
        RECT 198.000 -34.440 198.410 -34.000 ;
        RECT 201.180 -34.270 201.630 -33.990 ;
        RECT 205.000 -34.270 205.450 -33.990 ;
        RECT 214.680 -33.990 216.210 -33.780 ;
        RECT 216.590 -33.870 217.030 -33.780 ;
        RECT 199.010 -34.440 199.460 -34.360 ;
        RECT 197.160 -34.680 199.460 -34.440 ;
        RECT 197.160 -34.780 197.610 -34.680 ;
        RECT 199.010 -34.780 199.460 -34.680 ;
        RECT 200.410 -34.440 200.860 -34.330 ;
        RECT 202.260 -34.440 202.710 -34.330 ;
        RECT 200.410 -34.680 202.710 -34.440 ;
        RECT 200.410 -34.750 200.860 -34.680 ;
        RECT 183.660 -35.310 184.110 -35.260 ;
        RECT 182.020 -35.600 184.110 -35.310 ;
        RECT 182.020 -35.650 182.470 -35.600 ;
        RECT 165.270 -36.230 165.720 -36.160 ;
        RECT 163.420 -36.470 165.720 -36.230 ;
        RECT 163.420 -36.580 163.870 -36.470 ;
        RECT 165.270 -36.580 165.720 -36.470 ;
        RECT 166.670 -36.230 167.120 -36.130 ;
        RECT 168.520 -36.230 168.970 -36.130 ;
        RECT 166.670 -36.470 168.970 -36.230 ;
        RECT 166.670 -36.550 167.120 -36.470 ;
        RECT 147.180 -37.130 148.710 -36.920 ;
        RECT 149.090 -37.130 149.540 -37.040 ;
        RECT 149.920 -37.130 151.450 -36.920 ;
        RECT 160.680 -36.920 161.130 -36.640 ;
        RECT 164.500 -36.920 164.950 -36.640 ;
        RECT 167.720 -36.910 168.130 -36.470 ;
        RECT 168.520 -36.580 168.970 -36.470 ;
        RECT 170.160 -36.230 170.610 -36.130 ;
        RECT 172.010 -36.230 172.460 -36.130 ;
        RECT 170.160 -36.470 172.460 -36.230 ;
        RECT 170.160 -36.580 170.610 -36.470 ;
        RECT 171.000 -36.910 171.410 -36.470 ;
        RECT 172.010 -36.550 172.460 -36.470 ;
        RECT 173.410 -36.230 173.860 -36.160 ;
        RECT 174.460 -36.230 174.870 -35.800 ;
        RECT 175.260 -36.230 175.710 -36.130 ;
        RECT 173.410 -36.470 175.710 -36.230 ;
        RECT 173.410 -36.580 173.860 -36.470 ;
        RECT 175.260 -36.580 175.710 -36.470 ;
        RECT 176.920 -36.230 177.370 -36.130 ;
        RECT 177.760 -36.230 178.170 -35.800 ;
        RECT 180.920 -35.870 182.470 -35.650 ;
        RECT 182.850 -35.660 183.280 -35.600 ;
        RECT 183.660 -35.650 184.110 -35.600 ;
        RECT 184.710 -35.650 185.210 -35.260 ;
        RECT 183.660 -35.870 185.210 -35.650 ;
        RECT 194.420 -35.260 195.970 -35.040 ;
        RECT 194.420 -35.650 194.920 -35.260 ;
        RECT 195.520 -35.310 195.970 -35.260 ;
        RECT 196.350 -35.310 196.780 -35.250 ;
        RECT 197.160 -35.260 198.710 -35.040 ;
        RECT 201.460 -35.110 201.870 -34.680 ;
        RECT 202.260 -34.780 202.710 -34.680 ;
        RECT 203.920 -34.440 204.370 -34.330 ;
        RECT 205.770 -34.440 206.220 -34.330 ;
        RECT 203.920 -34.680 206.220 -34.440 ;
        RECT 203.920 -34.780 204.370 -34.680 ;
        RECT 204.760 -35.110 205.170 -34.680 ;
        RECT 205.770 -34.750 206.220 -34.680 ;
        RECT 207.170 -34.440 207.620 -34.360 ;
        RECT 208.220 -34.440 208.630 -34.000 ;
        RECT 209.020 -34.440 209.470 -34.330 ;
        RECT 207.170 -34.680 209.470 -34.440 ;
        RECT 207.170 -34.780 207.620 -34.680 ;
        RECT 209.020 -34.780 209.470 -34.680 ;
        RECT 210.660 -34.440 211.110 -34.330 ;
        RECT 211.500 -34.440 211.910 -34.000 ;
        RECT 214.680 -34.270 215.130 -33.990 ;
        RECT 212.510 -34.440 212.960 -34.360 ;
        RECT 210.660 -34.680 212.960 -34.440 ;
        RECT 210.660 -34.780 211.110 -34.680 ;
        RECT 212.510 -34.780 212.960 -34.680 ;
        RECT 213.910 -34.440 214.360 -34.330 ;
        RECT 215.760 -34.440 216.210 -34.330 ;
        RECT 213.910 -34.680 216.210 -34.440 ;
        RECT 213.910 -34.750 214.360 -34.680 ;
        RECT 197.160 -35.310 197.610 -35.260 ;
        RECT 195.520 -35.600 197.610 -35.310 ;
        RECT 195.520 -35.650 195.970 -35.600 ;
        RECT 178.770 -36.230 179.220 -36.160 ;
        RECT 176.920 -36.470 179.220 -36.230 ;
        RECT 176.920 -36.580 177.370 -36.470 ;
        RECT 178.770 -36.580 179.220 -36.470 ;
        RECT 180.170 -36.230 180.620 -36.130 ;
        RECT 182.020 -36.230 182.470 -36.130 ;
        RECT 180.170 -36.470 182.470 -36.230 ;
        RECT 180.170 -36.550 180.620 -36.470 ;
        RECT 160.680 -37.130 162.210 -36.920 ;
        RECT 162.590 -37.130 163.040 -37.040 ;
        RECT 163.420 -37.130 164.950 -36.920 ;
        RECT 174.180 -36.920 174.630 -36.640 ;
        RECT 178.000 -36.920 178.450 -36.640 ;
        RECT 181.220 -36.910 181.630 -36.470 ;
        RECT 182.020 -36.580 182.470 -36.470 ;
        RECT 183.660 -36.230 184.110 -36.130 ;
        RECT 185.510 -36.230 185.960 -36.130 ;
        RECT 183.660 -36.470 185.960 -36.230 ;
        RECT 183.660 -36.580 184.110 -36.470 ;
        RECT 184.500 -36.910 184.910 -36.470 ;
        RECT 185.510 -36.550 185.960 -36.470 ;
        RECT 186.910 -36.230 187.360 -36.160 ;
        RECT 187.960 -36.230 188.370 -35.800 ;
        RECT 188.760 -36.230 189.210 -36.130 ;
        RECT 186.910 -36.470 189.210 -36.230 ;
        RECT 186.910 -36.580 187.360 -36.470 ;
        RECT 188.760 -36.580 189.210 -36.470 ;
        RECT 190.420 -36.230 190.870 -36.130 ;
        RECT 191.260 -36.230 191.670 -35.800 ;
        RECT 194.420 -35.870 195.970 -35.650 ;
        RECT 196.350 -35.660 196.780 -35.600 ;
        RECT 197.160 -35.650 197.610 -35.600 ;
        RECT 198.210 -35.650 198.710 -35.260 ;
        RECT 197.160 -35.870 198.710 -35.650 ;
        RECT 207.920 -35.260 209.470 -35.040 ;
        RECT 207.920 -35.650 208.420 -35.260 ;
        RECT 209.020 -35.310 209.470 -35.260 ;
        RECT 209.850 -35.310 210.280 -35.250 ;
        RECT 210.660 -35.260 212.210 -35.040 ;
        RECT 214.960 -35.110 215.370 -34.680 ;
        RECT 215.760 -34.780 216.210 -34.680 ;
        RECT 210.660 -35.310 211.110 -35.260 ;
        RECT 209.020 -35.600 211.110 -35.310 ;
        RECT 209.020 -35.650 209.470 -35.600 ;
        RECT 192.270 -36.230 192.720 -36.160 ;
        RECT 190.420 -36.470 192.720 -36.230 ;
        RECT 190.420 -36.580 190.870 -36.470 ;
        RECT 192.270 -36.580 192.720 -36.470 ;
        RECT 193.670 -36.230 194.120 -36.130 ;
        RECT 195.520 -36.230 195.970 -36.130 ;
        RECT 193.670 -36.470 195.970 -36.230 ;
        RECT 193.670 -36.550 194.120 -36.470 ;
        RECT 174.180 -37.130 175.710 -36.920 ;
        RECT 176.090 -37.130 176.540 -37.040 ;
        RECT 176.920 -37.130 178.450 -36.920 ;
        RECT 187.680 -36.920 188.130 -36.640 ;
        RECT 191.500 -36.920 191.950 -36.640 ;
        RECT 194.720 -36.910 195.130 -36.470 ;
        RECT 195.520 -36.580 195.970 -36.470 ;
        RECT 197.160 -36.230 197.610 -36.130 ;
        RECT 199.010 -36.230 199.460 -36.130 ;
        RECT 197.160 -36.470 199.460 -36.230 ;
        RECT 197.160 -36.580 197.610 -36.470 ;
        RECT 198.000 -36.910 198.410 -36.470 ;
        RECT 199.010 -36.550 199.460 -36.470 ;
        RECT 200.410 -36.230 200.860 -36.160 ;
        RECT 201.460 -36.230 201.870 -35.800 ;
        RECT 202.260 -36.230 202.710 -36.130 ;
        RECT 200.410 -36.470 202.710 -36.230 ;
        RECT 200.410 -36.580 200.860 -36.470 ;
        RECT 202.260 -36.580 202.710 -36.470 ;
        RECT 203.920 -36.230 204.370 -36.130 ;
        RECT 204.760 -36.230 205.170 -35.800 ;
        RECT 207.920 -35.870 209.470 -35.650 ;
        RECT 209.850 -35.660 210.280 -35.600 ;
        RECT 210.660 -35.650 211.110 -35.600 ;
        RECT 211.710 -35.650 212.210 -35.260 ;
        RECT 210.660 -35.870 212.210 -35.650 ;
        RECT 205.770 -36.230 206.220 -36.160 ;
        RECT 203.920 -36.470 206.220 -36.230 ;
        RECT 203.920 -36.580 204.370 -36.470 ;
        RECT 205.770 -36.580 206.220 -36.470 ;
        RECT 207.170 -36.230 207.620 -36.130 ;
        RECT 209.020 -36.230 209.470 -36.130 ;
        RECT 207.170 -36.470 209.470 -36.230 ;
        RECT 207.170 -36.550 207.620 -36.470 ;
        RECT 187.680 -37.130 189.210 -36.920 ;
        RECT 189.590 -37.130 190.040 -37.040 ;
        RECT 190.420 -37.130 191.950 -36.920 ;
        RECT 201.180 -36.920 201.630 -36.640 ;
        RECT 205.000 -36.920 205.450 -36.640 ;
        RECT 208.220 -36.910 208.630 -36.470 ;
        RECT 209.020 -36.580 209.470 -36.470 ;
        RECT 210.660 -36.230 211.110 -36.130 ;
        RECT 212.510 -36.230 212.960 -36.130 ;
        RECT 210.660 -36.470 212.960 -36.230 ;
        RECT 210.660 -36.580 211.110 -36.470 ;
        RECT 211.500 -36.910 211.910 -36.470 ;
        RECT 212.510 -36.550 212.960 -36.470 ;
        RECT 213.910 -36.230 214.360 -36.160 ;
        RECT 214.960 -36.230 215.370 -35.800 ;
        RECT 215.760 -36.230 216.210 -36.130 ;
        RECT 213.910 -36.470 216.210 -36.230 ;
        RECT 213.910 -36.580 214.360 -36.470 ;
        RECT 215.760 -36.580 216.210 -36.470 ;
        RECT 201.180 -37.130 202.710 -36.920 ;
        RECT 203.090 -37.130 203.540 -37.040 ;
        RECT 203.920 -37.130 205.450 -36.920 ;
        RECT 214.680 -36.920 215.130 -36.640 ;
        RECT 214.680 -37.130 216.210 -36.920 ;
        RECT 216.590 -37.130 217.030 -37.040 ;
        RECT 13.260 -37.390 15.370 -37.130 ;
        RECT 26.760 -37.390 28.870 -37.130 ;
        RECT 40.260 -37.390 42.370 -37.130 ;
        RECT 53.760 -37.390 55.870 -37.130 ;
        RECT 67.260 -37.390 69.370 -37.130 ;
        RECT 80.760 -37.390 82.870 -37.130 ;
        RECT 94.260 -37.390 96.370 -37.130 ;
        RECT 107.760 -37.390 109.870 -37.130 ;
        RECT 121.260 -37.390 123.370 -37.130 ;
        RECT 134.760 -37.390 136.870 -37.130 ;
        RECT 148.260 -37.390 150.370 -37.130 ;
        RECT 161.760 -37.390 163.870 -37.130 ;
        RECT 175.260 -37.390 177.370 -37.130 ;
        RECT 188.760 -37.390 190.870 -37.130 ;
        RECT 202.260 -37.390 204.370 -37.130 ;
        RECT 215.760 -37.190 217.030 -37.130 ;
        RECT 215.760 -37.380 217.240 -37.190 ;
        RECT 215.760 -37.390 217.030 -37.380 ;
        RECT 12.180 -37.600 13.710 -37.390 ;
        RECT 14.090 -37.480 14.540 -37.390 ;
        RECT 14.920 -37.600 16.450 -37.390 ;
        RECT 1.420 -38.050 1.870 -37.940 ;
        RECT 3.270 -38.050 3.720 -37.940 ;
        RECT 1.420 -38.290 3.720 -38.050 ;
        RECT 1.420 -38.390 1.870 -38.290 ;
        RECT 2.260 -38.720 2.670 -38.290 ;
        RECT 3.270 -38.360 3.720 -38.290 ;
        RECT 4.670 -38.050 5.120 -37.970 ;
        RECT 5.720 -38.050 6.130 -37.610 ;
        RECT 6.520 -38.050 6.970 -37.940 ;
        RECT 4.670 -38.290 6.970 -38.050 ;
        RECT 4.670 -38.390 5.120 -38.290 ;
        RECT 6.520 -38.390 6.970 -38.290 ;
        RECT 8.160 -38.050 8.610 -37.940 ;
        RECT 9.000 -38.050 9.410 -37.610 ;
        RECT 12.180 -37.880 12.630 -37.600 ;
        RECT 16.000 -37.880 16.450 -37.600 ;
        RECT 25.680 -37.600 27.210 -37.390 ;
        RECT 27.590 -37.480 28.040 -37.390 ;
        RECT 28.420 -37.600 29.950 -37.390 ;
        RECT 10.010 -38.050 10.460 -37.970 ;
        RECT 8.160 -38.290 10.460 -38.050 ;
        RECT 8.160 -38.390 8.610 -38.290 ;
        RECT 10.010 -38.390 10.460 -38.290 ;
        RECT 11.410 -38.050 11.860 -37.940 ;
        RECT 13.260 -38.050 13.710 -37.940 ;
        RECT 11.410 -38.290 13.710 -38.050 ;
        RECT 11.410 -38.360 11.860 -38.290 ;
        RECT 5.420 -38.870 6.970 -38.650 ;
        RECT 5.420 -39.260 5.920 -38.870 ;
        RECT 6.520 -38.920 6.970 -38.870 ;
        RECT 7.350 -38.920 7.780 -38.860 ;
        RECT 8.160 -38.870 9.710 -38.650 ;
        RECT 12.460 -38.720 12.870 -38.290 ;
        RECT 13.260 -38.390 13.710 -38.290 ;
        RECT 14.920 -38.050 15.370 -37.940 ;
        RECT 16.770 -38.050 17.220 -37.940 ;
        RECT 14.920 -38.290 17.220 -38.050 ;
        RECT 14.920 -38.390 15.370 -38.290 ;
        RECT 15.760 -38.720 16.170 -38.290 ;
        RECT 16.770 -38.360 17.220 -38.290 ;
        RECT 18.170 -38.050 18.620 -37.970 ;
        RECT 19.220 -38.050 19.630 -37.610 ;
        RECT 20.020 -38.050 20.470 -37.940 ;
        RECT 18.170 -38.290 20.470 -38.050 ;
        RECT 18.170 -38.390 18.620 -38.290 ;
        RECT 20.020 -38.390 20.470 -38.290 ;
        RECT 21.660 -38.050 22.110 -37.940 ;
        RECT 22.500 -38.050 22.910 -37.610 ;
        RECT 25.680 -37.880 26.130 -37.600 ;
        RECT 29.500 -37.880 29.950 -37.600 ;
        RECT 39.180 -37.600 40.710 -37.390 ;
        RECT 41.090 -37.480 41.540 -37.390 ;
        RECT 41.920 -37.600 43.450 -37.390 ;
        RECT 23.510 -38.050 23.960 -37.970 ;
        RECT 21.660 -38.290 23.960 -38.050 ;
        RECT 21.660 -38.390 22.110 -38.290 ;
        RECT 23.510 -38.390 23.960 -38.290 ;
        RECT 24.910 -38.050 25.360 -37.940 ;
        RECT 26.760 -38.050 27.210 -37.940 ;
        RECT 24.910 -38.290 27.210 -38.050 ;
        RECT 24.910 -38.360 25.360 -38.290 ;
        RECT 8.160 -38.920 8.610 -38.870 ;
        RECT 6.520 -39.210 8.610 -38.920 ;
        RECT 6.520 -39.260 6.970 -39.210 ;
        RECT 1.420 -39.840 1.870 -39.740 ;
        RECT 2.260 -39.840 2.670 -39.410 ;
        RECT 5.420 -39.480 6.970 -39.260 ;
        RECT 7.350 -39.270 7.780 -39.210 ;
        RECT 8.160 -39.260 8.610 -39.210 ;
        RECT 9.210 -39.260 9.710 -38.870 ;
        RECT 8.160 -39.480 9.710 -39.260 ;
        RECT 18.920 -38.870 20.470 -38.650 ;
        RECT 18.920 -39.260 19.420 -38.870 ;
        RECT 20.020 -38.920 20.470 -38.870 ;
        RECT 20.850 -38.920 21.280 -38.860 ;
        RECT 21.660 -38.870 23.210 -38.650 ;
        RECT 25.960 -38.720 26.370 -38.290 ;
        RECT 26.760 -38.390 27.210 -38.290 ;
        RECT 28.420 -38.050 28.870 -37.940 ;
        RECT 30.270 -38.050 30.720 -37.940 ;
        RECT 28.420 -38.290 30.720 -38.050 ;
        RECT 28.420 -38.390 28.870 -38.290 ;
        RECT 29.260 -38.720 29.670 -38.290 ;
        RECT 30.270 -38.360 30.720 -38.290 ;
        RECT 31.670 -38.050 32.120 -37.970 ;
        RECT 32.720 -38.050 33.130 -37.610 ;
        RECT 33.520 -38.050 33.970 -37.940 ;
        RECT 31.670 -38.290 33.970 -38.050 ;
        RECT 31.670 -38.390 32.120 -38.290 ;
        RECT 33.520 -38.390 33.970 -38.290 ;
        RECT 35.160 -38.050 35.610 -37.940 ;
        RECT 36.000 -38.050 36.410 -37.610 ;
        RECT 39.180 -37.880 39.630 -37.600 ;
        RECT 43.000 -37.880 43.450 -37.600 ;
        RECT 52.680 -37.600 54.210 -37.390 ;
        RECT 54.590 -37.480 55.040 -37.390 ;
        RECT 55.420 -37.600 56.950 -37.390 ;
        RECT 37.010 -38.050 37.460 -37.970 ;
        RECT 35.160 -38.290 37.460 -38.050 ;
        RECT 35.160 -38.390 35.610 -38.290 ;
        RECT 37.010 -38.390 37.460 -38.290 ;
        RECT 38.410 -38.050 38.860 -37.940 ;
        RECT 40.260 -38.050 40.710 -37.940 ;
        RECT 38.410 -38.290 40.710 -38.050 ;
        RECT 38.410 -38.360 38.860 -38.290 ;
        RECT 21.660 -38.920 22.110 -38.870 ;
        RECT 20.020 -39.210 22.110 -38.920 ;
        RECT 20.020 -39.260 20.470 -39.210 ;
        RECT 3.270 -39.840 3.720 -39.770 ;
        RECT 1.420 -40.080 3.720 -39.840 ;
        RECT 1.420 -40.190 1.870 -40.080 ;
        RECT 3.270 -40.190 3.720 -40.080 ;
        RECT 4.670 -39.840 5.120 -39.740 ;
        RECT 6.520 -39.840 6.970 -39.740 ;
        RECT 4.670 -40.080 6.970 -39.840 ;
        RECT 4.670 -40.160 5.120 -40.080 ;
        RECT 5.720 -40.520 6.130 -40.080 ;
        RECT 6.520 -40.190 6.970 -40.080 ;
        RECT 8.160 -39.840 8.610 -39.740 ;
        RECT 10.010 -39.840 10.460 -39.740 ;
        RECT 8.160 -40.080 10.460 -39.840 ;
        RECT 8.160 -40.190 8.610 -40.080 ;
        RECT 9.000 -40.520 9.410 -40.080 ;
        RECT 10.010 -40.160 10.460 -40.080 ;
        RECT 11.410 -39.840 11.860 -39.770 ;
        RECT 12.460 -39.840 12.870 -39.410 ;
        RECT 13.260 -39.840 13.710 -39.740 ;
        RECT 11.410 -40.080 13.710 -39.840 ;
        RECT 11.410 -40.190 11.860 -40.080 ;
        RECT 13.260 -40.190 13.710 -40.080 ;
        RECT 14.920 -39.840 15.370 -39.740 ;
        RECT 15.760 -39.840 16.170 -39.410 ;
        RECT 18.920 -39.480 20.470 -39.260 ;
        RECT 20.850 -39.270 21.280 -39.210 ;
        RECT 21.660 -39.260 22.110 -39.210 ;
        RECT 22.710 -39.260 23.210 -38.870 ;
        RECT 21.660 -39.480 23.210 -39.260 ;
        RECT 32.420 -38.870 33.970 -38.650 ;
        RECT 32.420 -39.260 32.920 -38.870 ;
        RECT 33.520 -38.920 33.970 -38.870 ;
        RECT 34.350 -38.920 34.780 -38.860 ;
        RECT 35.160 -38.870 36.710 -38.650 ;
        RECT 39.460 -38.720 39.870 -38.290 ;
        RECT 40.260 -38.390 40.710 -38.290 ;
        RECT 41.920 -38.050 42.370 -37.940 ;
        RECT 43.770 -38.050 44.220 -37.940 ;
        RECT 41.920 -38.290 44.220 -38.050 ;
        RECT 41.920 -38.390 42.370 -38.290 ;
        RECT 42.760 -38.720 43.170 -38.290 ;
        RECT 43.770 -38.360 44.220 -38.290 ;
        RECT 45.170 -38.050 45.620 -37.970 ;
        RECT 46.220 -38.050 46.630 -37.610 ;
        RECT 47.020 -38.050 47.470 -37.940 ;
        RECT 45.170 -38.290 47.470 -38.050 ;
        RECT 45.170 -38.390 45.620 -38.290 ;
        RECT 47.020 -38.390 47.470 -38.290 ;
        RECT 48.660 -38.050 49.110 -37.940 ;
        RECT 49.500 -38.050 49.910 -37.610 ;
        RECT 52.680 -37.880 53.130 -37.600 ;
        RECT 56.500 -37.880 56.950 -37.600 ;
        RECT 66.180 -37.600 67.710 -37.390 ;
        RECT 68.090 -37.480 68.540 -37.390 ;
        RECT 68.920 -37.600 70.450 -37.390 ;
        RECT 50.510 -38.050 50.960 -37.970 ;
        RECT 48.660 -38.290 50.960 -38.050 ;
        RECT 48.660 -38.390 49.110 -38.290 ;
        RECT 50.510 -38.390 50.960 -38.290 ;
        RECT 51.910 -38.050 52.360 -37.940 ;
        RECT 53.760 -38.050 54.210 -37.940 ;
        RECT 51.910 -38.290 54.210 -38.050 ;
        RECT 51.910 -38.360 52.360 -38.290 ;
        RECT 35.160 -38.920 35.610 -38.870 ;
        RECT 33.520 -39.210 35.610 -38.920 ;
        RECT 33.520 -39.260 33.970 -39.210 ;
        RECT 16.770 -39.840 17.220 -39.770 ;
        RECT 14.920 -40.080 17.220 -39.840 ;
        RECT 14.920 -40.190 15.370 -40.080 ;
        RECT 16.770 -40.190 17.220 -40.080 ;
        RECT 18.170 -39.840 18.620 -39.740 ;
        RECT 20.020 -39.840 20.470 -39.740 ;
        RECT 18.170 -40.080 20.470 -39.840 ;
        RECT 18.170 -40.160 18.620 -40.080 ;
        RECT 12.180 -40.530 12.630 -40.250 ;
        RECT 16.000 -40.530 16.450 -40.250 ;
        RECT 19.220 -40.520 19.630 -40.080 ;
        RECT 20.020 -40.190 20.470 -40.080 ;
        RECT 21.660 -39.840 22.110 -39.740 ;
        RECT 23.510 -39.840 23.960 -39.740 ;
        RECT 21.660 -40.080 23.960 -39.840 ;
        RECT 21.660 -40.190 22.110 -40.080 ;
        RECT 22.500 -40.520 22.910 -40.080 ;
        RECT 23.510 -40.160 23.960 -40.080 ;
        RECT 24.910 -39.840 25.360 -39.770 ;
        RECT 25.960 -39.840 26.370 -39.410 ;
        RECT 26.760 -39.840 27.210 -39.740 ;
        RECT 24.910 -40.080 27.210 -39.840 ;
        RECT 24.910 -40.190 25.360 -40.080 ;
        RECT 26.760 -40.190 27.210 -40.080 ;
        RECT 28.420 -39.840 28.870 -39.740 ;
        RECT 29.260 -39.840 29.670 -39.410 ;
        RECT 32.420 -39.480 33.970 -39.260 ;
        RECT 34.350 -39.270 34.780 -39.210 ;
        RECT 35.160 -39.260 35.610 -39.210 ;
        RECT 36.210 -39.260 36.710 -38.870 ;
        RECT 35.160 -39.480 36.710 -39.260 ;
        RECT 45.920 -38.870 47.470 -38.650 ;
        RECT 45.920 -39.260 46.420 -38.870 ;
        RECT 47.020 -38.920 47.470 -38.870 ;
        RECT 47.850 -38.920 48.280 -38.860 ;
        RECT 48.660 -38.870 50.210 -38.650 ;
        RECT 52.960 -38.720 53.370 -38.290 ;
        RECT 53.760 -38.390 54.210 -38.290 ;
        RECT 55.420 -38.050 55.870 -37.940 ;
        RECT 57.270 -38.050 57.720 -37.940 ;
        RECT 55.420 -38.290 57.720 -38.050 ;
        RECT 55.420 -38.390 55.870 -38.290 ;
        RECT 56.260 -38.720 56.670 -38.290 ;
        RECT 57.270 -38.360 57.720 -38.290 ;
        RECT 58.670 -38.050 59.120 -37.970 ;
        RECT 59.720 -38.050 60.130 -37.610 ;
        RECT 60.520 -38.050 60.970 -37.940 ;
        RECT 58.670 -38.290 60.970 -38.050 ;
        RECT 58.670 -38.390 59.120 -38.290 ;
        RECT 60.520 -38.390 60.970 -38.290 ;
        RECT 62.160 -38.050 62.610 -37.940 ;
        RECT 63.000 -38.050 63.410 -37.610 ;
        RECT 66.180 -37.880 66.630 -37.600 ;
        RECT 70.000 -37.880 70.450 -37.600 ;
        RECT 79.680 -37.600 81.210 -37.390 ;
        RECT 81.590 -37.480 82.040 -37.390 ;
        RECT 82.420 -37.600 83.950 -37.390 ;
        RECT 64.010 -38.050 64.460 -37.970 ;
        RECT 62.160 -38.290 64.460 -38.050 ;
        RECT 62.160 -38.390 62.610 -38.290 ;
        RECT 64.010 -38.390 64.460 -38.290 ;
        RECT 65.410 -38.050 65.860 -37.940 ;
        RECT 67.260 -38.050 67.710 -37.940 ;
        RECT 65.410 -38.290 67.710 -38.050 ;
        RECT 65.410 -38.360 65.860 -38.290 ;
        RECT 48.660 -38.920 49.110 -38.870 ;
        RECT 47.020 -39.210 49.110 -38.920 ;
        RECT 47.020 -39.260 47.470 -39.210 ;
        RECT 30.270 -39.840 30.720 -39.770 ;
        RECT 28.420 -40.080 30.720 -39.840 ;
        RECT 28.420 -40.190 28.870 -40.080 ;
        RECT 30.270 -40.190 30.720 -40.080 ;
        RECT 31.670 -39.840 32.120 -39.740 ;
        RECT 33.520 -39.840 33.970 -39.740 ;
        RECT 31.670 -40.080 33.970 -39.840 ;
        RECT 31.670 -40.160 32.120 -40.080 ;
        RECT 12.180 -40.740 13.710 -40.530 ;
        RECT 13.260 -40.750 13.710 -40.740 ;
        RECT 14.090 -40.750 14.540 -40.660 ;
        RECT 14.920 -40.740 16.450 -40.530 ;
        RECT 25.680 -40.530 26.130 -40.250 ;
        RECT 29.500 -40.530 29.950 -40.250 ;
        RECT 32.720 -40.520 33.130 -40.080 ;
        RECT 33.520 -40.190 33.970 -40.080 ;
        RECT 35.160 -39.840 35.610 -39.740 ;
        RECT 37.010 -39.840 37.460 -39.740 ;
        RECT 35.160 -40.080 37.460 -39.840 ;
        RECT 35.160 -40.190 35.610 -40.080 ;
        RECT 36.000 -40.520 36.410 -40.080 ;
        RECT 37.010 -40.160 37.460 -40.080 ;
        RECT 38.410 -39.840 38.860 -39.770 ;
        RECT 39.460 -39.840 39.870 -39.410 ;
        RECT 40.260 -39.840 40.710 -39.740 ;
        RECT 38.410 -40.080 40.710 -39.840 ;
        RECT 38.410 -40.190 38.860 -40.080 ;
        RECT 40.260 -40.190 40.710 -40.080 ;
        RECT 41.920 -39.840 42.370 -39.740 ;
        RECT 42.760 -39.840 43.170 -39.410 ;
        RECT 45.920 -39.480 47.470 -39.260 ;
        RECT 47.850 -39.270 48.280 -39.210 ;
        RECT 48.660 -39.260 49.110 -39.210 ;
        RECT 49.710 -39.260 50.210 -38.870 ;
        RECT 48.660 -39.480 50.210 -39.260 ;
        RECT 59.420 -38.870 60.970 -38.650 ;
        RECT 59.420 -39.260 59.920 -38.870 ;
        RECT 60.520 -38.920 60.970 -38.870 ;
        RECT 61.350 -38.920 61.780 -38.860 ;
        RECT 62.160 -38.870 63.710 -38.650 ;
        RECT 66.460 -38.720 66.870 -38.290 ;
        RECT 67.260 -38.390 67.710 -38.290 ;
        RECT 68.920 -38.050 69.370 -37.940 ;
        RECT 70.770 -38.050 71.220 -37.940 ;
        RECT 68.920 -38.290 71.220 -38.050 ;
        RECT 68.920 -38.390 69.370 -38.290 ;
        RECT 69.760 -38.720 70.170 -38.290 ;
        RECT 70.770 -38.360 71.220 -38.290 ;
        RECT 72.170 -38.050 72.620 -37.970 ;
        RECT 73.220 -38.050 73.630 -37.610 ;
        RECT 74.020 -38.050 74.470 -37.940 ;
        RECT 72.170 -38.290 74.470 -38.050 ;
        RECT 72.170 -38.390 72.620 -38.290 ;
        RECT 74.020 -38.390 74.470 -38.290 ;
        RECT 75.660 -38.050 76.110 -37.940 ;
        RECT 76.500 -38.050 76.910 -37.610 ;
        RECT 79.680 -37.880 80.130 -37.600 ;
        RECT 83.500 -37.880 83.950 -37.600 ;
        RECT 93.180 -37.600 94.710 -37.390 ;
        RECT 95.090 -37.480 95.540 -37.390 ;
        RECT 95.920 -37.600 97.450 -37.390 ;
        RECT 77.510 -38.050 77.960 -37.970 ;
        RECT 75.660 -38.290 77.960 -38.050 ;
        RECT 75.660 -38.390 76.110 -38.290 ;
        RECT 77.510 -38.390 77.960 -38.290 ;
        RECT 78.910 -38.050 79.360 -37.940 ;
        RECT 80.760 -38.050 81.210 -37.940 ;
        RECT 78.910 -38.290 81.210 -38.050 ;
        RECT 78.910 -38.360 79.360 -38.290 ;
        RECT 62.160 -38.920 62.610 -38.870 ;
        RECT 60.520 -39.210 62.610 -38.920 ;
        RECT 60.520 -39.260 60.970 -39.210 ;
        RECT 43.770 -39.840 44.220 -39.770 ;
        RECT 41.920 -40.080 44.220 -39.840 ;
        RECT 41.920 -40.190 42.370 -40.080 ;
        RECT 43.770 -40.190 44.220 -40.080 ;
        RECT 45.170 -39.840 45.620 -39.740 ;
        RECT 47.020 -39.840 47.470 -39.740 ;
        RECT 45.170 -40.080 47.470 -39.840 ;
        RECT 45.170 -40.160 45.620 -40.080 ;
        RECT 25.680 -40.740 27.210 -40.530 ;
        RECT 14.920 -40.750 15.370 -40.740 ;
        RECT 13.260 -41.000 15.370 -40.750 ;
        RECT 13.260 -41.100 13.710 -41.000 ;
        RECT 14.090 -41.090 14.540 -41.000 ;
        RECT 14.920 -41.100 15.370 -41.000 ;
        RECT 26.760 -40.750 27.210 -40.740 ;
        RECT 27.590 -40.750 28.040 -40.660 ;
        RECT 28.420 -40.740 29.950 -40.530 ;
        RECT 39.180 -40.530 39.630 -40.250 ;
        RECT 43.000 -40.530 43.450 -40.250 ;
        RECT 46.220 -40.520 46.630 -40.080 ;
        RECT 47.020 -40.190 47.470 -40.080 ;
        RECT 48.660 -39.840 49.110 -39.740 ;
        RECT 50.510 -39.840 50.960 -39.740 ;
        RECT 48.660 -40.080 50.960 -39.840 ;
        RECT 48.660 -40.190 49.110 -40.080 ;
        RECT 49.500 -40.520 49.910 -40.080 ;
        RECT 50.510 -40.160 50.960 -40.080 ;
        RECT 51.910 -39.840 52.360 -39.770 ;
        RECT 52.960 -39.840 53.370 -39.410 ;
        RECT 53.760 -39.840 54.210 -39.740 ;
        RECT 51.910 -40.080 54.210 -39.840 ;
        RECT 51.910 -40.190 52.360 -40.080 ;
        RECT 53.760 -40.190 54.210 -40.080 ;
        RECT 55.420 -39.840 55.870 -39.740 ;
        RECT 56.260 -39.840 56.670 -39.410 ;
        RECT 59.420 -39.480 60.970 -39.260 ;
        RECT 61.350 -39.270 61.780 -39.210 ;
        RECT 62.160 -39.260 62.610 -39.210 ;
        RECT 63.210 -39.260 63.710 -38.870 ;
        RECT 62.160 -39.480 63.710 -39.260 ;
        RECT 72.920 -38.870 74.470 -38.650 ;
        RECT 72.920 -39.260 73.420 -38.870 ;
        RECT 74.020 -38.920 74.470 -38.870 ;
        RECT 74.850 -38.920 75.280 -38.860 ;
        RECT 75.660 -38.870 77.210 -38.650 ;
        RECT 79.960 -38.720 80.370 -38.290 ;
        RECT 80.760 -38.390 81.210 -38.290 ;
        RECT 82.420 -38.050 82.870 -37.940 ;
        RECT 84.270 -38.050 84.720 -37.940 ;
        RECT 82.420 -38.290 84.720 -38.050 ;
        RECT 82.420 -38.390 82.870 -38.290 ;
        RECT 83.260 -38.720 83.670 -38.290 ;
        RECT 84.270 -38.360 84.720 -38.290 ;
        RECT 85.670 -38.050 86.120 -37.970 ;
        RECT 86.720 -38.050 87.130 -37.610 ;
        RECT 87.520 -38.050 87.970 -37.940 ;
        RECT 85.670 -38.290 87.970 -38.050 ;
        RECT 85.670 -38.390 86.120 -38.290 ;
        RECT 87.520 -38.390 87.970 -38.290 ;
        RECT 89.160 -38.050 89.610 -37.940 ;
        RECT 90.000 -38.050 90.410 -37.610 ;
        RECT 93.180 -37.880 93.630 -37.600 ;
        RECT 97.000 -37.880 97.450 -37.600 ;
        RECT 106.680 -37.600 108.210 -37.390 ;
        RECT 108.590 -37.480 109.040 -37.390 ;
        RECT 109.420 -37.600 110.950 -37.390 ;
        RECT 91.010 -38.050 91.460 -37.970 ;
        RECT 89.160 -38.290 91.460 -38.050 ;
        RECT 89.160 -38.390 89.610 -38.290 ;
        RECT 91.010 -38.390 91.460 -38.290 ;
        RECT 92.410 -38.050 92.860 -37.940 ;
        RECT 94.260 -38.050 94.710 -37.940 ;
        RECT 92.410 -38.290 94.710 -38.050 ;
        RECT 92.410 -38.360 92.860 -38.290 ;
        RECT 75.660 -38.920 76.110 -38.870 ;
        RECT 74.020 -39.210 76.110 -38.920 ;
        RECT 74.020 -39.260 74.470 -39.210 ;
        RECT 57.270 -39.840 57.720 -39.770 ;
        RECT 55.420 -40.080 57.720 -39.840 ;
        RECT 55.420 -40.190 55.870 -40.080 ;
        RECT 57.270 -40.190 57.720 -40.080 ;
        RECT 58.670 -39.840 59.120 -39.740 ;
        RECT 60.520 -39.840 60.970 -39.740 ;
        RECT 58.670 -40.080 60.970 -39.840 ;
        RECT 58.670 -40.160 59.120 -40.080 ;
        RECT 39.180 -40.740 40.710 -40.530 ;
        RECT 28.420 -40.750 28.870 -40.740 ;
        RECT 26.760 -41.000 28.870 -40.750 ;
        RECT 26.760 -41.100 27.210 -41.000 ;
        RECT 27.590 -41.090 28.040 -41.000 ;
        RECT 28.420 -41.100 28.870 -41.000 ;
        RECT 40.260 -40.750 40.710 -40.740 ;
        RECT 41.090 -40.750 41.540 -40.660 ;
        RECT 41.920 -40.740 43.450 -40.530 ;
        RECT 52.680 -40.530 53.130 -40.250 ;
        RECT 56.500 -40.530 56.950 -40.250 ;
        RECT 59.720 -40.520 60.130 -40.080 ;
        RECT 60.520 -40.190 60.970 -40.080 ;
        RECT 62.160 -39.840 62.610 -39.740 ;
        RECT 64.010 -39.840 64.460 -39.740 ;
        RECT 62.160 -40.080 64.460 -39.840 ;
        RECT 62.160 -40.190 62.610 -40.080 ;
        RECT 63.000 -40.520 63.410 -40.080 ;
        RECT 64.010 -40.160 64.460 -40.080 ;
        RECT 65.410 -39.840 65.860 -39.770 ;
        RECT 66.460 -39.840 66.870 -39.410 ;
        RECT 67.260 -39.840 67.710 -39.740 ;
        RECT 65.410 -40.080 67.710 -39.840 ;
        RECT 65.410 -40.190 65.860 -40.080 ;
        RECT 67.260 -40.190 67.710 -40.080 ;
        RECT 68.920 -39.840 69.370 -39.740 ;
        RECT 69.760 -39.840 70.170 -39.410 ;
        RECT 72.920 -39.480 74.470 -39.260 ;
        RECT 74.850 -39.270 75.280 -39.210 ;
        RECT 75.660 -39.260 76.110 -39.210 ;
        RECT 76.710 -39.260 77.210 -38.870 ;
        RECT 75.660 -39.480 77.210 -39.260 ;
        RECT 86.420 -38.870 87.970 -38.650 ;
        RECT 86.420 -39.260 86.920 -38.870 ;
        RECT 87.520 -38.920 87.970 -38.870 ;
        RECT 88.350 -38.920 88.780 -38.860 ;
        RECT 89.160 -38.870 90.710 -38.650 ;
        RECT 93.460 -38.720 93.870 -38.290 ;
        RECT 94.260 -38.390 94.710 -38.290 ;
        RECT 95.920 -38.050 96.370 -37.940 ;
        RECT 97.770 -38.050 98.220 -37.940 ;
        RECT 95.920 -38.290 98.220 -38.050 ;
        RECT 95.920 -38.390 96.370 -38.290 ;
        RECT 96.760 -38.720 97.170 -38.290 ;
        RECT 97.770 -38.360 98.220 -38.290 ;
        RECT 99.170 -38.050 99.620 -37.970 ;
        RECT 100.220 -38.050 100.630 -37.610 ;
        RECT 101.020 -38.050 101.470 -37.940 ;
        RECT 99.170 -38.290 101.470 -38.050 ;
        RECT 99.170 -38.390 99.620 -38.290 ;
        RECT 101.020 -38.390 101.470 -38.290 ;
        RECT 102.660 -38.050 103.110 -37.940 ;
        RECT 103.500 -38.050 103.910 -37.610 ;
        RECT 106.680 -37.880 107.130 -37.600 ;
        RECT 110.500 -37.880 110.950 -37.600 ;
        RECT 120.180 -37.600 121.710 -37.390 ;
        RECT 122.090 -37.480 122.540 -37.390 ;
        RECT 122.920 -37.600 124.450 -37.390 ;
        RECT 104.510 -38.050 104.960 -37.970 ;
        RECT 102.660 -38.290 104.960 -38.050 ;
        RECT 102.660 -38.390 103.110 -38.290 ;
        RECT 104.510 -38.390 104.960 -38.290 ;
        RECT 105.910 -38.050 106.360 -37.940 ;
        RECT 107.760 -38.050 108.210 -37.940 ;
        RECT 105.910 -38.290 108.210 -38.050 ;
        RECT 105.910 -38.360 106.360 -38.290 ;
        RECT 89.160 -38.920 89.610 -38.870 ;
        RECT 87.520 -39.210 89.610 -38.920 ;
        RECT 87.520 -39.260 87.970 -39.210 ;
        RECT 70.770 -39.840 71.220 -39.770 ;
        RECT 68.920 -40.080 71.220 -39.840 ;
        RECT 68.920 -40.190 69.370 -40.080 ;
        RECT 70.770 -40.190 71.220 -40.080 ;
        RECT 72.170 -39.840 72.620 -39.740 ;
        RECT 74.020 -39.840 74.470 -39.740 ;
        RECT 72.170 -40.080 74.470 -39.840 ;
        RECT 72.170 -40.160 72.620 -40.080 ;
        RECT 52.680 -40.730 54.210 -40.530 ;
        RECT 54.590 -40.730 55.040 -40.660 ;
        RECT 55.420 -40.730 56.950 -40.530 ;
        RECT 52.680 -40.740 56.950 -40.730 ;
        RECT 66.180 -40.530 66.630 -40.250 ;
        RECT 70.000 -40.530 70.450 -40.250 ;
        RECT 73.220 -40.520 73.630 -40.080 ;
        RECT 74.020 -40.190 74.470 -40.080 ;
        RECT 75.660 -39.840 76.110 -39.740 ;
        RECT 77.510 -39.840 77.960 -39.740 ;
        RECT 75.660 -40.080 77.960 -39.840 ;
        RECT 75.660 -40.190 76.110 -40.080 ;
        RECT 76.500 -40.520 76.910 -40.080 ;
        RECT 77.510 -40.160 77.960 -40.080 ;
        RECT 78.910 -39.840 79.360 -39.770 ;
        RECT 79.960 -39.840 80.370 -39.410 ;
        RECT 80.760 -39.840 81.210 -39.740 ;
        RECT 78.910 -40.080 81.210 -39.840 ;
        RECT 78.910 -40.190 79.360 -40.080 ;
        RECT 80.760 -40.190 81.210 -40.080 ;
        RECT 82.420 -39.840 82.870 -39.740 ;
        RECT 83.260 -39.840 83.670 -39.410 ;
        RECT 86.420 -39.480 87.970 -39.260 ;
        RECT 88.350 -39.270 88.780 -39.210 ;
        RECT 89.160 -39.260 89.610 -39.210 ;
        RECT 90.210 -39.260 90.710 -38.870 ;
        RECT 89.160 -39.480 90.710 -39.260 ;
        RECT 99.920 -38.870 101.470 -38.650 ;
        RECT 99.920 -39.260 100.420 -38.870 ;
        RECT 101.020 -38.920 101.470 -38.870 ;
        RECT 101.850 -38.920 102.280 -38.860 ;
        RECT 102.660 -38.870 104.210 -38.650 ;
        RECT 106.960 -38.720 107.370 -38.290 ;
        RECT 107.760 -38.390 108.210 -38.290 ;
        RECT 109.420 -38.050 109.870 -37.940 ;
        RECT 111.270 -38.050 111.720 -37.940 ;
        RECT 109.420 -38.290 111.720 -38.050 ;
        RECT 109.420 -38.390 109.870 -38.290 ;
        RECT 110.260 -38.720 110.670 -38.290 ;
        RECT 111.270 -38.360 111.720 -38.290 ;
        RECT 112.670 -38.050 113.120 -37.970 ;
        RECT 113.720 -38.050 114.130 -37.610 ;
        RECT 114.520 -38.050 114.970 -37.940 ;
        RECT 112.670 -38.290 114.970 -38.050 ;
        RECT 112.670 -38.390 113.120 -38.290 ;
        RECT 114.520 -38.390 114.970 -38.290 ;
        RECT 116.160 -38.050 116.610 -37.940 ;
        RECT 117.000 -38.050 117.410 -37.610 ;
        RECT 120.180 -37.880 120.630 -37.600 ;
        RECT 124.000 -37.880 124.450 -37.600 ;
        RECT 133.680 -37.600 135.210 -37.390 ;
        RECT 135.590 -37.480 136.040 -37.390 ;
        RECT 136.420 -37.600 137.950 -37.390 ;
        RECT 118.010 -38.050 118.460 -37.970 ;
        RECT 116.160 -38.290 118.460 -38.050 ;
        RECT 116.160 -38.390 116.610 -38.290 ;
        RECT 118.010 -38.390 118.460 -38.290 ;
        RECT 119.410 -38.050 119.860 -37.940 ;
        RECT 121.260 -38.050 121.710 -37.940 ;
        RECT 119.410 -38.290 121.710 -38.050 ;
        RECT 119.410 -38.360 119.860 -38.290 ;
        RECT 102.660 -38.920 103.110 -38.870 ;
        RECT 101.020 -39.210 103.110 -38.920 ;
        RECT 101.020 -39.260 101.470 -39.210 ;
        RECT 84.270 -39.840 84.720 -39.770 ;
        RECT 82.420 -40.080 84.720 -39.840 ;
        RECT 82.420 -40.190 82.870 -40.080 ;
        RECT 84.270 -40.190 84.720 -40.080 ;
        RECT 85.670 -39.840 86.120 -39.740 ;
        RECT 87.520 -39.840 87.970 -39.740 ;
        RECT 85.670 -40.080 87.970 -39.840 ;
        RECT 85.670 -40.160 86.120 -40.080 ;
        RECT 66.180 -40.740 67.710 -40.530 ;
        RECT 41.920 -40.750 42.370 -40.740 ;
        RECT 40.260 -41.000 42.370 -40.750 ;
        RECT 40.260 -41.100 40.710 -41.000 ;
        RECT 41.090 -41.090 41.540 -41.000 ;
        RECT 41.920 -41.100 42.370 -41.000 ;
        RECT 53.760 -41.050 55.870 -40.740 ;
        RECT 53.760 -41.100 54.210 -41.050 ;
        RECT 54.590 -41.090 55.040 -41.050 ;
        RECT 55.420 -41.100 55.870 -41.050 ;
        RECT 67.260 -40.750 67.710 -40.740 ;
        RECT 68.090 -40.750 68.540 -40.660 ;
        RECT 68.920 -40.740 70.450 -40.530 ;
        RECT 79.680 -40.530 80.130 -40.250 ;
        RECT 83.500 -40.530 83.950 -40.250 ;
        RECT 86.720 -40.520 87.130 -40.080 ;
        RECT 87.520 -40.190 87.970 -40.080 ;
        RECT 89.160 -39.840 89.610 -39.740 ;
        RECT 91.010 -39.840 91.460 -39.740 ;
        RECT 89.160 -40.080 91.460 -39.840 ;
        RECT 89.160 -40.190 89.610 -40.080 ;
        RECT 90.000 -40.520 90.410 -40.080 ;
        RECT 91.010 -40.160 91.460 -40.080 ;
        RECT 92.410 -39.840 92.860 -39.770 ;
        RECT 93.460 -39.840 93.870 -39.410 ;
        RECT 94.260 -39.840 94.710 -39.740 ;
        RECT 92.410 -40.080 94.710 -39.840 ;
        RECT 92.410 -40.190 92.860 -40.080 ;
        RECT 94.260 -40.190 94.710 -40.080 ;
        RECT 95.920 -39.840 96.370 -39.740 ;
        RECT 96.760 -39.840 97.170 -39.410 ;
        RECT 99.920 -39.480 101.470 -39.260 ;
        RECT 101.850 -39.270 102.280 -39.210 ;
        RECT 102.660 -39.260 103.110 -39.210 ;
        RECT 103.710 -39.260 104.210 -38.870 ;
        RECT 102.660 -39.480 104.210 -39.260 ;
        RECT 113.420 -38.870 114.970 -38.650 ;
        RECT 113.420 -39.260 113.920 -38.870 ;
        RECT 114.520 -38.920 114.970 -38.870 ;
        RECT 115.350 -38.920 115.780 -38.860 ;
        RECT 116.160 -38.870 117.710 -38.650 ;
        RECT 120.460 -38.720 120.870 -38.290 ;
        RECT 121.260 -38.390 121.710 -38.290 ;
        RECT 122.920 -38.050 123.370 -37.940 ;
        RECT 124.770 -38.050 125.220 -37.940 ;
        RECT 122.920 -38.290 125.220 -38.050 ;
        RECT 122.920 -38.390 123.370 -38.290 ;
        RECT 123.760 -38.720 124.170 -38.290 ;
        RECT 124.770 -38.360 125.220 -38.290 ;
        RECT 126.170 -38.050 126.620 -37.970 ;
        RECT 127.220 -38.050 127.630 -37.610 ;
        RECT 128.020 -38.050 128.470 -37.940 ;
        RECT 126.170 -38.290 128.470 -38.050 ;
        RECT 126.170 -38.390 126.620 -38.290 ;
        RECT 128.020 -38.390 128.470 -38.290 ;
        RECT 129.660 -38.050 130.110 -37.940 ;
        RECT 130.500 -38.050 130.910 -37.610 ;
        RECT 133.680 -37.880 134.130 -37.600 ;
        RECT 137.500 -37.880 137.950 -37.600 ;
        RECT 147.180 -37.600 148.710 -37.390 ;
        RECT 149.090 -37.480 149.540 -37.390 ;
        RECT 149.920 -37.600 151.450 -37.390 ;
        RECT 131.510 -38.050 131.960 -37.970 ;
        RECT 129.660 -38.290 131.960 -38.050 ;
        RECT 129.660 -38.390 130.110 -38.290 ;
        RECT 131.510 -38.390 131.960 -38.290 ;
        RECT 132.910 -38.050 133.360 -37.940 ;
        RECT 134.760 -38.050 135.210 -37.940 ;
        RECT 132.910 -38.290 135.210 -38.050 ;
        RECT 132.910 -38.360 133.360 -38.290 ;
        RECT 116.160 -38.920 116.610 -38.870 ;
        RECT 114.520 -39.210 116.610 -38.920 ;
        RECT 114.520 -39.260 114.970 -39.210 ;
        RECT 97.770 -39.840 98.220 -39.770 ;
        RECT 95.920 -40.080 98.220 -39.840 ;
        RECT 95.920 -40.190 96.370 -40.080 ;
        RECT 97.770 -40.190 98.220 -40.080 ;
        RECT 99.170 -39.840 99.620 -39.740 ;
        RECT 101.020 -39.840 101.470 -39.740 ;
        RECT 99.170 -40.080 101.470 -39.840 ;
        RECT 99.170 -40.160 99.620 -40.080 ;
        RECT 79.680 -40.740 81.210 -40.530 ;
        RECT 68.920 -40.750 69.370 -40.740 ;
        RECT 67.260 -41.000 69.370 -40.750 ;
        RECT 67.260 -41.100 67.710 -41.000 ;
        RECT 68.090 -41.090 68.540 -41.000 ;
        RECT 68.920 -41.100 69.370 -41.000 ;
        RECT 80.760 -40.750 81.210 -40.740 ;
        RECT 81.590 -40.750 82.040 -40.660 ;
        RECT 82.420 -40.740 83.950 -40.530 ;
        RECT 93.180 -40.530 93.630 -40.250 ;
        RECT 97.000 -40.530 97.450 -40.250 ;
        RECT 100.220 -40.520 100.630 -40.080 ;
        RECT 101.020 -40.190 101.470 -40.080 ;
        RECT 102.660 -39.840 103.110 -39.740 ;
        RECT 104.510 -39.840 104.960 -39.740 ;
        RECT 102.660 -40.080 104.960 -39.840 ;
        RECT 102.660 -40.190 103.110 -40.080 ;
        RECT 103.500 -40.520 103.910 -40.080 ;
        RECT 104.510 -40.160 104.960 -40.080 ;
        RECT 105.910 -39.840 106.360 -39.770 ;
        RECT 106.960 -39.840 107.370 -39.410 ;
        RECT 107.760 -39.840 108.210 -39.740 ;
        RECT 105.910 -40.080 108.210 -39.840 ;
        RECT 105.910 -40.190 106.360 -40.080 ;
        RECT 107.760 -40.190 108.210 -40.080 ;
        RECT 109.420 -39.840 109.870 -39.740 ;
        RECT 110.260 -39.840 110.670 -39.410 ;
        RECT 113.420 -39.480 114.970 -39.260 ;
        RECT 115.350 -39.270 115.780 -39.210 ;
        RECT 116.160 -39.260 116.610 -39.210 ;
        RECT 117.210 -39.260 117.710 -38.870 ;
        RECT 116.160 -39.480 117.710 -39.260 ;
        RECT 126.920 -38.870 128.470 -38.650 ;
        RECT 126.920 -39.260 127.420 -38.870 ;
        RECT 128.020 -38.920 128.470 -38.870 ;
        RECT 128.850 -38.920 129.280 -38.860 ;
        RECT 129.660 -38.870 131.210 -38.650 ;
        RECT 133.960 -38.720 134.370 -38.290 ;
        RECT 134.760 -38.390 135.210 -38.290 ;
        RECT 136.420 -38.050 136.870 -37.940 ;
        RECT 138.270 -38.050 138.720 -37.940 ;
        RECT 136.420 -38.290 138.720 -38.050 ;
        RECT 136.420 -38.390 136.870 -38.290 ;
        RECT 137.260 -38.720 137.670 -38.290 ;
        RECT 138.270 -38.360 138.720 -38.290 ;
        RECT 139.670 -38.050 140.120 -37.970 ;
        RECT 140.720 -38.050 141.130 -37.610 ;
        RECT 141.520 -38.050 141.970 -37.940 ;
        RECT 139.670 -38.290 141.970 -38.050 ;
        RECT 139.670 -38.390 140.120 -38.290 ;
        RECT 141.520 -38.390 141.970 -38.290 ;
        RECT 143.160 -38.050 143.610 -37.940 ;
        RECT 144.000 -38.050 144.410 -37.610 ;
        RECT 147.180 -37.880 147.630 -37.600 ;
        RECT 151.000 -37.880 151.450 -37.600 ;
        RECT 160.680 -37.600 162.210 -37.390 ;
        RECT 162.590 -37.480 163.040 -37.390 ;
        RECT 163.420 -37.600 164.950 -37.390 ;
        RECT 145.010 -38.050 145.460 -37.970 ;
        RECT 143.160 -38.290 145.460 -38.050 ;
        RECT 143.160 -38.390 143.610 -38.290 ;
        RECT 145.010 -38.390 145.460 -38.290 ;
        RECT 146.410 -38.050 146.860 -37.940 ;
        RECT 148.260 -38.050 148.710 -37.940 ;
        RECT 146.410 -38.290 148.710 -38.050 ;
        RECT 146.410 -38.360 146.860 -38.290 ;
        RECT 129.660 -38.920 130.110 -38.870 ;
        RECT 128.020 -39.210 130.110 -38.920 ;
        RECT 128.020 -39.260 128.470 -39.210 ;
        RECT 111.270 -39.840 111.720 -39.770 ;
        RECT 109.420 -40.080 111.720 -39.840 ;
        RECT 109.420 -40.190 109.870 -40.080 ;
        RECT 111.270 -40.190 111.720 -40.080 ;
        RECT 112.670 -39.840 113.120 -39.740 ;
        RECT 114.520 -39.840 114.970 -39.740 ;
        RECT 112.670 -40.080 114.970 -39.840 ;
        RECT 112.670 -40.160 113.120 -40.080 ;
        RECT 93.180 -40.740 94.710 -40.530 ;
        RECT 82.420 -40.750 82.870 -40.740 ;
        RECT 80.760 -41.000 82.870 -40.750 ;
        RECT 80.760 -41.100 81.210 -41.000 ;
        RECT 81.590 -41.090 82.040 -41.000 ;
        RECT 82.420 -41.100 82.870 -41.000 ;
        RECT 94.260 -40.750 94.710 -40.740 ;
        RECT 95.090 -40.750 95.540 -40.660 ;
        RECT 95.920 -40.740 97.450 -40.530 ;
        RECT 106.680 -40.530 107.130 -40.250 ;
        RECT 110.500 -40.530 110.950 -40.250 ;
        RECT 113.720 -40.520 114.130 -40.080 ;
        RECT 114.520 -40.190 114.970 -40.080 ;
        RECT 116.160 -39.840 116.610 -39.740 ;
        RECT 118.010 -39.840 118.460 -39.740 ;
        RECT 116.160 -40.080 118.460 -39.840 ;
        RECT 116.160 -40.190 116.610 -40.080 ;
        RECT 117.000 -40.520 117.410 -40.080 ;
        RECT 118.010 -40.160 118.460 -40.080 ;
        RECT 119.410 -39.840 119.860 -39.770 ;
        RECT 120.460 -39.840 120.870 -39.410 ;
        RECT 121.260 -39.840 121.710 -39.740 ;
        RECT 119.410 -40.080 121.710 -39.840 ;
        RECT 119.410 -40.190 119.860 -40.080 ;
        RECT 121.260 -40.190 121.710 -40.080 ;
        RECT 122.920 -39.840 123.370 -39.740 ;
        RECT 123.760 -39.840 124.170 -39.410 ;
        RECT 126.920 -39.480 128.470 -39.260 ;
        RECT 128.850 -39.270 129.280 -39.210 ;
        RECT 129.660 -39.260 130.110 -39.210 ;
        RECT 130.710 -39.260 131.210 -38.870 ;
        RECT 129.660 -39.480 131.210 -39.260 ;
        RECT 140.420 -38.870 141.970 -38.650 ;
        RECT 140.420 -39.260 140.920 -38.870 ;
        RECT 141.520 -38.920 141.970 -38.870 ;
        RECT 142.350 -38.920 142.780 -38.860 ;
        RECT 143.160 -38.870 144.710 -38.650 ;
        RECT 147.460 -38.720 147.870 -38.290 ;
        RECT 148.260 -38.390 148.710 -38.290 ;
        RECT 149.920 -38.050 150.370 -37.940 ;
        RECT 151.770 -38.050 152.220 -37.940 ;
        RECT 149.920 -38.290 152.220 -38.050 ;
        RECT 149.920 -38.390 150.370 -38.290 ;
        RECT 150.760 -38.720 151.170 -38.290 ;
        RECT 151.770 -38.360 152.220 -38.290 ;
        RECT 153.170 -38.050 153.620 -37.970 ;
        RECT 154.220 -38.050 154.630 -37.610 ;
        RECT 155.020 -38.050 155.470 -37.940 ;
        RECT 153.170 -38.290 155.470 -38.050 ;
        RECT 153.170 -38.390 153.620 -38.290 ;
        RECT 155.020 -38.390 155.470 -38.290 ;
        RECT 156.660 -38.050 157.110 -37.940 ;
        RECT 157.500 -38.050 157.910 -37.610 ;
        RECT 160.680 -37.880 161.130 -37.600 ;
        RECT 164.500 -37.880 164.950 -37.600 ;
        RECT 174.180 -37.600 175.710 -37.390 ;
        RECT 176.090 -37.480 176.540 -37.390 ;
        RECT 176.920 -37.600 178.450 -37.390 ;
        RECT 158.510 -38.050 158.960 -37.970 ;
        RECT 156.660 -38.290 158.960 -38.050 ;
        RECT 156.660 -38.390 157.110 -38.290 ;
        RECT 158.510 -38.390 158.960 -38.290 ;
        RECT 159.910 -38.050 160.360 -37.940 ;
        RECT 161.760 -38.050 162.210 -37.940 ;
        RECT 159.910 -38.290 162.210 -38.050 ;
        RECT 159.910 -38.360 160.360 -38.290 ;
        RECT 143.160 -38.920 143.610 -38.870 ;
        RECT 141.520 -39.210 143.610 -38.920 ;
        RECT 141.520 -39.260 141.970 -39.210 ;
        RECT 124.770 -39.840 125.220 -39.770 ;
        RECT 122.920 -40.080 125.220 -39.840 ;
        RECT 122.920 -40.190 123.370 -40.080 ;
        RECT 124.770 -40.190 125.220 -40.080 ;
        RECT 126.170 -39.840 126.620 -39.740 ;
        RECT 128.020 -39.840 128.470 -39.740 ;
        RECT 126.170 -40.080 128.470 -39.840 ;
        RECT 126.170 -40.160 126.620 -40.080 ;
        RECT 106.680 -40.730 108.210 -40.530 ;
        RECT 108.590 -40.730 109.040 -40.660 ;
        RECT 109.420 -40.730 110.950 -40.530 ;
        RECT 106.680 -40.740 110.950 -40.730 ;
        RECT 120.180 -40.530 120.630 -40.250 ;
        RECT 124.000 -40.530 124.450 -40.250 ;
        RECT 127.220 -40.520 127.630 -40.080 ;
        RECT 128.020 -40.190 128.470 -40.080 ;
        RECT 129.660 -39.840 130.110 -39.740 ;
        RECT 131.510 -39.840 131.960 -39.740 ;
        RECT 129.660 -40.080 131.960 -39.840 ;
        RECT 129.660 -40.190 130.110 -40.080 ;
        RECT 130.500 -40.520 130.910 -40.080 ;
        RECT 131.510 -40.160 131.960 -40.080 ;
        RECT 132.910 -39.840 133.360 -39.770 ;
        RECT 133.960 -39.840 134.370 -39.410 ;
        RECT 134.760 -39.840 135.210 -39.740 ;
        RECT 132.910 -40.080 135.210 -39.840 ;
        RECT 132.910 -40.190 133.360 -40.080 ;
        RECT 134.760 -40.190 135.210 -40.080 ;
        RECT 136.420 -39.840 136.870 -39.740 ;
        RECT 137.260 -39.840 137.670 -39.410 ;
        RECT 140.420 -39.480 141.970 -39.260 ;
        RECT 142.350 -39.270 142.780 -39.210 ;
        RECT 143.160 -39.260 143.610 -39.210 ;
        RECT 144.210 -39.260 144.710 -38.870 ;
        RECT 143.160 -39.480 144.710 -39.260 ;
        RECT 153.920 -38.870 155.470 -38.650 ;
        RECT 153.920 -39.260 154.420 -38.870 ;
        RECT 155.020 -38.920 155.470 -38.870 ;
        RECT 155.850 -38.920 156.280 -38.860 ;
        RECT 156.660 -38.870 158.210 -38.650 ;
        RECT 160.960 -38.720 161.370 -38.290 ;
        RECT 161.760 -38.390 162.210 -38.290 ;
        RECT 163.420 -38.050 163.870 -37.940 ;
        RECT 165.270 -38.050 165.720 -37.940 ;
        RECT 163.420 -38.290 165.720 -38.050 ;
        RECT 163.420 -38.390 163.870 -38.290 ;
        RECT 164.260 -38.720 164.670 -38.290 ;
        RECT 165.270 -38.360 165.720 -38.290 ;
        RECT 166.670 -38.050 167.120 -37.970 ;
        RECT 167.720 -38.050 168.130 -37.610 ;
        RECT 168.520 -38.050 168.970 -37.940 ;
        RECT 166.670 -38.290 168.970 -38.050 ;
        RECT 166.670 -38.390 167.120 -38.290 ;
        RECT 168.520 -38.390 168.970 -38.290 ;
        RECT 170.160 -38.050 170.610 -37.940 ;
        RECT 171.000 -38.050 171.410 -37.610 ;
        RECT 174.180 -37.880 174.630 -37.600 ;
        RECT 178.000 -37.880 178.450 -37.600 ;
        RECT 187.680 -37.600 189.210 -37.390 ;
        RECT 189.590 -37.480 190.040 -37.390 ;
        RECT 190.420 -37.600 191.950 -37.390 ;
        RECT 172.010 -38.050 172.460 -37.970 ;
        RECT 170.160 -38.290 172.460 -38.050 ;
        RECT 170.160 -38.390 170.610 -38.290 ;
        RECT 172.010 -38.390 172.460 -38.290 ;
        RECT 173.410 -38.050 173.860 -37.940 ;
        RECT 175.260 -38.050 175.710 -37.940 ;
        RECT 173.410 -38.290 175.710 -38.050 ;
        RECT 173.410 -38.360 173.860 -38.290 ;
        RECT 156.660 -38.920 157.110 -38.870 ;
        RECT 155.020 -39.210 157.110 -38.920 ;
        RECT 155.020 -39.260 155.470 -39.210 ;
        RECT 138.270 -39.840 138.720 -39.770 ;
        RECT 136.420 -40.080 138.720 -39.840 ;
        RECT 136.420 -40.190 136.870 -40.080 ;
        RECT 138.270 -40.190 138.720 -40.080 ;
        RECT 139.670 -39.840 140.120 -39.740 ;
        RECT 141.520 -39.840 141.970 -39.740 ;
        RECT 139.670 -40.080 141.970 -39.840 ;
        RECT 139.670 -40.160 140.120 -40.080 ;
        RECT 120.180 -40.740 121.710 -40.530 ;
        RECT 95.920 -40.750 96.370 -40.740 ;
        RECT 94.260 -41.000 96.370 -40.750 ;
        RECT 94.260 -41.100 94.710 -41.000 ;
        RECT 95.090 -41.090 95.540 -41.000 ;
        RECT 95.920 -41.100 96.370 -41.000 ;
        RECT 107.760 -41.050 109.870 -40.740 ;
        RECT 107.760 -41.100 108.210 -41.050 ;
        RECT 108.590 -41.090 109.040 -41.050 ;
        RECT 109.420 -41.100 109.870 -41.050 ;
        RECT 121.260 -40.750 121.710 -40.740 ;
        RECT 122.090 -40.750 122.540 -40.660 ;
        RECT 122.920 -40.740 124.450 -40.530 ;
        RECT 133.680 -40.530 134.130 -40.250 ;
        RECT 137.500 -40.530 137.950 -40.250 ;
        RECT 140.720 -40.520 141.130 -40.080 ;
        RECT 141.520 -40.190 141.970 -40.080 ;
        RECT 143.160 -39.840 143.610 -39.740 ;
        RECT 145.010 -39.840 145.460 -39.740 ;
        RECT 143.160 -40.080 145.460 -39.840 ;
        RECT 143.160 -40.190 143.610 -40.080 ;
        RECT 144.000 -40.520 144.410 -40.080 ;
        RECT 145.010 -40.160 145.460 -40.080 ;
        RECT 146.410 -39.840 146.860 -39.770 ;
        RECT 147.460 -39.840 147.870 -39.410 ;
        RECT 148.260 -39.840 148.710 -39.740 ;
        RECT 146.410 -40.080 148.710 -39.840 ;
        RECT 146.410 -40.190 146.860 -40.080 ;
        RECT 148.260 -40.190 148.710 -40.080 ;
        RECT 149.920 -39.840 150.370 -39.740 ;
        RECT 150.760 -39.840 151.170 -39.410 ;
        RECT 153.920 -39.480 155.470 -39.260 ;
        RECT 155.850 -39.270 156.280 -39.210 ;
        RECT 156.660 -39.260 157.110 -39.210 ;
        RECT 157.710 -39.260 158.210 -38.870 ;
        RECT 156.660 -39.480 158.210 -39.260 ;
        RECT 167.420 -38.870 168.970 -38.650 ;
        RECT 167.420 -39.260 167.920 -38.870 ;
        RECT 168.520 -38.920 168.970 -38.870 ;
        RECT 169.350 -38.920 169.780 -38.860 ;
        RECT 170.160 -38.870 171.710 -38.650 ;
        RECT 174.460 -38.720 174.870 -38.290 ;
        RECT 175.260 -38.390 175.710 -38.290 ;
        RECT 176.920 -38.050 177.370 -37.940 ;
        RECT 178.770 -38.050 179.220 -37.940 ;
        RECT 176.920 -38.290 179.220 -38.050 ;
        RECT 176.920 -38.390 177.370 -38.290 ;
        RECT 177.760 -38.720 178.170 -38.290 ;
        RECT 178.770 -38.360 179.220 -38.290 ;
        RECT 180.170 -38.050 180.620 -37.970 ;
        RECT 181.220 -38.050 181.630 -37.610 ;
        RECT 182.020 -38.050 182.470 -37.940 ;
        RECT 180.170 -38.290 182.470 -38.050 ;
        RECT 180.170 -38.390 180.620 -38.290 ;
        RECT 182.020 -38.390 182.470 -38.290 ;
        RECT 183.660 -38.050 184.110 -37.940 ;
        RECT 184.500 -38.050 184.910 -37.610 ;
        RECT 187.680 -37.880 188.130 -37.600 ;
        RECT 191.500 -37.880 191.950 -37.600 ;
        RECT 201.180 -37.600 202.710 -37.390 ;
        RECT 203.090 -37.480 203.540 -37.390 ;
        RECT 203.920 -37.600 205.450 -37.390 ;
        RECT 185.510 -38.050 185.960 -37.970 ;
        RECT 183.660 -38.290 185.960 -38.050 ;
        RECT 183.660 -38.390 184.110 -38.290 ;
        RECT 185.510 -38.390 185.960 -38.290 ;
        RECT 186.910 -38.050 187.360 -37.940 ;
        RECT 188.760 -38.050 189.210 -37.940 ;
        RECT 186.910 -38.290 189.210 -38.050 ;
        RECT 186.910 -38.360 187.360 -38.290 ;
        RECT 170.160 -38.920 170.610 -38.870 ;
        RECT 168.520 -39.210 170.610 -38.920 ;
        RECT 168.520 -39.260 168.970 -39.210 ;
        RECT 151.770 -39.840 152.220 -39.770 ;
        RECT 149.920 -40.080 152.220 -39.840 ;
        RECT 149.920 -40.190 150.370 -40.080 ;
        RECT 151.770 -40.190 152.220 -40.080 ;
        RECT 153.170 -39.840 153.620 -39.740 ;
        RECT 155.020 -39.840 155.470 -39.740 ;
        RECT 153.170 -40.080 155.470 -39.840 ;
        RECT 153.170 -40.160 153.620 -40.080 ;
        RECT 133.680 -40.740 135.210 -40.530 ;
        RECT 122.920 -40.750 123.370 -40.740 ;
        RECT 121.260 -41.000 123.370 -40.750 ;
        RECT 121.260 -41.100 121.710 -41.000 ;
        RECT 122.090 -41.090 122.540 -41.000 ;
        RECT 122.920 -41.100 123.370 -41.000 ;
        RECT 134.760 -40.750 135.210 -40.740 ;
        RECT 135.590 -40.750 136.040 -40.660 ;
        RECT 136.420 -40.740 137.950 -40.530 ;
        RECT 147.180 -40.530 147.630 -40.250 ;
        RECT 151.000 -40.530 151.450 -40.250 ;
        RECT 154.220 -40.520 154.630 -40.080 ;
        RECT 155.020 -40.190 155.470 -40.080 ;
        RECT 156.660 -39.840 157.110 -39.740 ;
        RECT 158.510 -39.840 158.960 -39.740 ;
        RECT 156.660 -40.080 158.960 -39.840 ;
        RECT 156.660 -40.190 157.110 -40.080 ;
        RECT 157.500 -40.520 157.910 -40.080 ;
        RECT 158.510 -40.160 158.960 -40.080 ;
        RECT 159.910 -39.840 160.360 -39.770 ;
        RECT 160.960 -39.840 161.370 -39.410 ;
        RECT 161.760 -39.840 162.210 -39.740 ;
        RECT 159.910 -40.080 162.210 -39.840 ;
        RECT 159.910 -40.190 160.360 -40.080 ;
        RECT 161.760 -40.190 162.210 -40.080 ;
        RECT 163.420 -39.840 163.870 -39.740 ;
        RECT 164.260 -39.840 164.670 -39.410 ;
        RECT 167.420 -39.480 168.970 -39.260 ;
        RECT 169.350 -39.270 169.780 -39.210 ;
        RECT 170.160 -39.260 170.610 -39.210 ;
        RECT 171.210 -39.260 171.710 -38.870 ;
        RECT 170.160 -39.480 171.710 -39.260 ;
        RECT 180.920 -38.870 182.470 -38.650 ;
        RECT 180.920 -39.260 181.420 -38.870 ;
        RECT 182.020 -38.920 182.470 -38.870 ;
        RECT 182.850 -38.920 183.280 -38.860 ;
        RECT 183.660 -38.870 185.210 -38.650 ;
        RECT 187.960 -38.720 188.370 -38.290 ;
        RECT 188.760 -38.390 189.210 -38.290 ;
        RECT 190.420 -38.050 190.870 -37.940 ;
        RECT 192.270 -38.050 192.720 -37.940 ;
        RECT 190.420 -38.290 192.720 -38.050 ;
        RECT 190.420 -38.390 190.870 -38.290 ;
        RECT 191.260 -38.720 191.670 -38.290 ;
        RECT 192.270 -38.360 192.720 -38.290 ;
        RECT 193.670 -38.050 194.120 -37.970 ;
        RECT 194.720 -38.050 195.130 -37.610 ;
        RECT 195.520 -38.050 195.970 -37.940 ;
        RECT 193.670 -38.290 195.970 -38.050 ;
        RECT 193.670 -38.390 194.120 -38.290 ;
        RECT 195.520 -38.390 195.970 -38.290 ;
        RECT 197.160 -38.050 197.610 -37.940 ;
        RECT 198.000 -38.050 198.410 -37.610 ;
        RECT 201.180 -37.880 201.630 -37.600 ;
        RECT 205.000 -37.880 205.450 -37.600 ;
        RECT 214.680 -37.600 216.210 -37.390 ;
        RECT 216.590 -37.480 217.030 -37.390 ;
        RECT 199.010 -38.050 199.460 -37.970 ;
        RECT 197.160 -38.290 199.460 -38.050 ;
        RECT 197.160 -38.390 197.610 -38.290 ;
        RECT 199.010 -38.390 199.460 -38.290 ;
        RECT 200.410 -38.050 200.860 -37.940 ;
        RECT 202.260 -38.050 202.710 -37.940 ;
        RECT 200.410 -38.290 202.710 -38.050 ;
        RECT 200.410 -38.360 200.860 -38.290 ;
        RECT 183.660 -38.920 184.110 -38.870 ;
        RECT 182.020 -39.210 184.110 -38.920 ;
        RECT 182.020 -39.260 182.470 -39.210 ;
        RECT 165.270 -39.840 165.720 -39.770 ;
        RECT 163.420 -40.080 165.720 -39.840 ;
        RECT 163.420 -40.190 163.870 -40.080 ;
        RECT 165.270 -40.190 165.720 -40.080 ;
        RECT 166.670 -39.840 167.120 -39.740 ;
        RECT 168.520 -39.840 168.970 -39.740 ;
        RECT 166.670 -40.080 168.970 -39.840 ;
        RECT 166.670 -40.160 167.120 -40.080 ;
        RECT 147.180 -40.740 148.710 -40.530 ;
        RECT 136.420 -40.750 136.870 -40.740 ;
        RECT 134.760 -41.000 136.870 -40.750 ;
        RECT 134.760 -41.100 135.210 -41.000 ;
        RECT 135.590 -41.090 136.040 -41.000 ;
        RECT 136.420 -41.100 136.870 -41.000 ;
        RECT 148.260 -40.750 148.710 -40.740 ;
        RECT 149.090 -40.750 149.540 -40.660 ;
        RECT 149.920 -40.740 151.450 -40.530 ;
        RECT 160.680 -40.530 161.130 -40.250 ;
        RECT 164.500 -40.530 164.950 -40.250 ;
        RECT 167.720 -40.520 168.130 -40.080 ;
        RECT 168.520 -40.190 168.970 -40.080 ;
        RECT 170.160 -39.840 170.610 -39.740 ;
        RECT 172.010 -39.840 172.460 -39.740 ;
        RECT 170.160 -40.080 172.460 -39.840 ;
        RECT 170.160 -40.190 170.610 -40.080 ;
        RECT 171.000 -40.520 171.410 -40.080 ;
        RECT 172.010 -40.160 172.460 -40.080 ;
        RECT 173.410 -39.840 173.860 -39.770 ;
        RECT 174.460 -39.840 174.870 -39.410 ;
        RECT 175.260 -39.840 175.710 -39.740 ;
        RECT 173.410 -40.080 175.710 -39.840 ;
        RECT 173.410 -40.190 173.860 -40.080 ;
        RECT 175.260 -40.190 175.710 -40.080 ;
        RECT 176.920 -39.840 177.370 -39.740 ;
        RECT 177.760 -39.840 178.170 -39.410 ;
        RECT 180.920 -39.480 182.470 -39.260 ;
        RECT 182.850 -39.270 183.280 -39.210 ;
        RECT 183.660 -39.260 184.110 -39.210 ;
        RECT 184.710 -39.260 185.210 -38.870 ;
        RECT 183.660 -39.480 185.210 -39.260 ;
        RECT 194.420 -38.870 195.970 -38.650 ;
        RECT 194.420 -39.260 194.920 -38.870 ;
        RECT 195.520 -38.920 195.970 -38.870 ;
        RECT 196.350 -38.920 196.780 -38.860 ;
        RECT 197.160 -38.870 198.710 -38.650 ;
        RECT 201.460 -38.720 201.870 -38.290 ;
        RECT 202.260 -38.390 202.710 -38.290 ;
        RECT 203.920 -38.050 204.370 -37.940 ;
        RECT 205.770 -38.050 206.220 -37.940 ;
        RECT 203.920 -38.290 206.220 -38.050 ;
        RECT 203.920 -38.390 204.370 -38.290 ;
        RECT 204.760 -38.720 205.170 -38.290 ;
        RECT 205.770 -38.360 206.220 -38.290 ;
        RECT 207.170 -38.050 207.620 -37.970 ;
        RECT 208.220 -38.050 208.630 -37.610 ;
        RECT 209.020 -38.050 209.470 -37.940 ;
        RECT 207.170 -38.290 209.470 -38.050 ;
        RECT 207.170 -38.390 207.620 -38.290 ;
        RECT 209.020 -38.390 209.470 -38.290 ;
        RECT 210.660 -38.050 211.110 -37.940 ;
        RECT 211.500 -38.050 211.910 -37.610 ;
        RECT 214.680 -37.880 215.130 -37.600 ;
        RECT 212.510 -38.050 212.960 -37.970 ;
        RECT 210.660 -38.290 212.960 -38.050 ;
        RECT 210.660 -38.390 211.110 -38.290 ;
        RECT 212.510 -38.390 212.960 -38.290 ;
        RECT 213.910 -38.050 214.360 -37.940 ;
        RECT 215.760 -38.050 216.210 -37.940 ;
        RECT 213.910 -38.290 216.210 -38.050 ;
        RECT 213.910 -38.360 214.360 -38.290 ;
        RECT 197.160 -38.920 197.610 -38.870 ;
        RECT 195.520 -39.210 197.610 -38.920 ;
        RECT 195.520 -39.260 195.970 -39.210 ;
        RECT 178.770 -39.840 179.220 -39.770 ;
        RECT 176.920 -40.080 179.220 -39.840 ;
        RECT 176.920 -40.190 177.370 -40.080 ;
        RECT 178.770 -40.190 179.220 -40.080 ;
        RECT 180.170 -39.840 180.620 -39.740 ;
        RECT 182.020 -39.840 182.470 -39.740 ;
        RECT 180.170 -40.080 182.470 -39.840 ;
        RECT 180.170 -40.160 180.620 -40.080 ;
        RECT 160.680 -40.730 162.210 -40.530 ;
        RECT 162.590 -40.730 163.040 -40.660 ;
        RECT 163.420 -40.730 164.950 -40.530 ;
        RECT 160.680 -40.740 164.950 -40.730 ;
        RECT 174.180 -40.530 174.630 -40.250 ;
        RECT 178.000 -40.530 178.450 -40.250 ;
        RECT 181.220 -40.520 181.630 -40.080 ;
        RECT 182.020 -40.190 182.470 -40.080 ;
        RECT 183.660 -39.840 184.110 -39.740 ;
        RECT 185.510 -39.840 185.960 -39.740 ;
        RECT 183.660 -40.080 185.960 -39.840 ;
        RECT 183.660 -40.190 184.110 -40.080 ;
        RECT 184.500 -40.520 184.910 -40.080 ;
        RECT 185.510 -40.160 185.960 -40.080 ;
        RECT 186.910 -39.840 187.360 -39.770 ;
        RECT 187.960 -39.840 188.370 -39.410 ;
        RECT 188.760 -39.840 189.210 -39.740 ;
        RECT 186.910 -40.080 189.210 -39.840 ;
        RECT 186.910 -40.190 187.360 -40.080 ;
        RECT 188.760 -40.190 189.210 -40.080 ;
        RECT 190.420 -39.840 190.870 -39.740 ;
        RECT 191.260 -39.840 191.670 -39.410 ;
        RECT 194.420 -39.480 195.970 -39.260 ;
        RECT 196.350 -39.270 196.780 -39.210 ;
        RECT 197.160 -39.260 197.610 -39.210 ;
        RECT 198.210 -39.260 198.710 -38.870 ;
        RECT 197.160 -39.480 198.710 -39.260 ;
        RECT 207.920 -38.870 209.470 -38.650 ;
        RECT 207.920 -39.260 208.420 -38.870 ;
        RECT 209.020 -38.920 209.470 -38.870 ;
        RECT 209.850 -38.920 210.280 -38.860 ;
        RECT 210.660 -38.870 212.210 -38.650 ;
        RECT 214.960 -38.720 215.370 -38.290 ;
        RECT 215.760 -38.390 216.210 -38.290 ;
        RECT 210.660 -38.920 211.110 -38.870 ;
        RECT 209.020 -39.210 211.110 -38.920 ;
        RECT 209.020 -39.260 209.470 -39.210 ;
        RECT 192.270 -39.840 192.720 -39.770 ;
        RECT 190.420 -40.080 192.720 -39.840 ;
        RECT 190.420 -40.190 190.870 -40.080 ;
        RECT 192.270 -40.190 192.720 -40.080 ;
        RECT 193.670 -39.840 194.120 -39.740 ;
        RECT 195.520 -39.840 195.970 -39.740 ;
        RECT 193.670 -40.080 195.970 -39.840 ;
        RECT 193.670 -40.160 194.120 -40.080 ;
        RECT 174.180 -40.740 175.710 -40.530 ;
        RECT 149.920 -40.750 150.370 -40.740 ;
        RECT 148.260 -41.000 150.370 -40.750 ;
        RECT 148.260 -41.100 148.710 -41.000 ;
        RECT 149.090 -41.090 149.540 -41.000 ;
        RECT 149.920 -41.100 150.370 -41.000 ;
        RECT 161.760 -41.050 163.870 -40.740 ;
        RECT 161.760 -41.100 162.210 -41.050 ;
        RECT 162.590 -41.090 163.040 -41.050 ;
        RECT 163.420 -41.100 163.870 -41.050 ;
        RECT 175.260 -40.750 175.710 -40.740 ;
        RECT 176.090 -40.750 176.540 -40.660 ;
        RECT 176.920 -40.740 178.450 -40.530 ;
        RECT 187.680 -40.530 188.130 -40.250 ;
        RECT 191.500 -40.530 191.950 -40.250 ;
        RECT 194.720 -40.520 195.130 -40.080 ;
        RECT 195.520 -40.190 195.970 -40.080 ;
        RECT 197.160 -39.840 197.610 -39.740 ;
        RECT 199.010 -39.840 199.460 -39.740 ;
        RECT 197.160 -40.080 199.460 -39.840 ;
        RECT 197.160 -40.190 197.610 -40.080 ;
        RECT 198.000 -40.520 198.410 -40.080 ;
        RECT 199.010 -40.160 199.460 -40.080 ;
        RECT 200.410 -39.840 200.860 -39.770 ;
        RECT 201.460 -39.840 201.870 -39.410 ;
        RECT 202.260 -39.840 202.710 -39.740 ;
        RECT 200.410 -40.080 202.710 -39.840 ;
        RECT 200.410 -40.190 200.860 -40.080 ;
        RECT 202.260 -40.190 202.710 -40.080 ;
        RECT 203.920 -39.840 204.370 -39.740 ;
        RECT 204.760 -39.840 205.170 -39.410 ;
        RECT 207.920 -39.480 209.470 -39.260 ;
        RECT 209.850 -39.270 210.280 -39.210 ;
        RECT 210.660 -39.260 211.110 -39.210 ;
        RECT 211.710 -39.260 212.210 -38.870 ;
        RECT 210.660 -39.480 212.210 -39.260 ;
        RECT 205.770 -39.840 206.220 -39.770 ;
        RECT 203.920 -40.080 206.220 -39.840 ;
        RECT 203.920 -40.190 204.370 -40.080 ;
        RECT 205.770 -40.190 206.220 -40.080 ;
        RECT 207.170 -39.840 207.620 -39.740 ;
        RECT 209.020 -39.840 209.470 -39.740 ;
        RECT 207.170 -40.080 209.470 -39.840 ;
        RECT 207.170 -40.160 207.620 -40.080 ;
        RECT 187.680 -40.740 189.210 -40.530 ;
        RECT 176.920 -40.750 177.370 -40.740 ;
        RECT 175.260 -41.000 177.370 -40.750 ;
        RECT 175.260 -41.100 175.710 -41.000 ;
        RECT 176.090 -41.090 176.540 -41.000 ;
        RECT 176.920 -41.100 177.370 -41.000 ;
        RECT 188.760 -40.750 189.210 -40.740 ;
        RECT 189.590 -40.750 190.040 -40.660 ;
        RECT 190.420 -40.740 191.950 -40.530 ;
        RECT 201.180 -40.530 201.630 -40.250 ;
        RECT 205.000 -40.530 205.450 -40.250 ;
        RECT 208.220 -40.520 208.630 -40.080 ;
        RECT 209.020 -40.190 209.470 -40.080 ;
        RECT 210.660 -39.840 211.110 -39.740 ;
        RECT 212.510 -39.840 212.960 -39.740 ;
        RECT 210.660 -40.080 212.960 -39.840 ;
        RECT 210.660 -40.190 211.110 -40.080 ;
        RECT 211.500 -40.520 211.910 -40.080 ;
        RECT 212.510 -40.160 212.960 -40.080 ;
        RECT 213.910 -39.840 214.360 -39.770 ;
        RECT 214.960 -39.840 215.370 -39.410 ;
        RECT 215.760 -39.840 216.210 -39.740 ;
        RECT 213.910 -40.080 216.210 -39.840 ;
        RECT 213.910 -40.190 214.360 -40.080 ;
        RECT 215.760 -40.190 216.210 -40.080 ;
        RECT 201.180 -40.740 202.710 -40.530 ;
        RECT 190.420 -40.750 190.870 -40.740 ;
        RECT 188.760 -41.000 190.870 -40.750 ;
        RECT 188.760 -41.100 189.210 -41.000 ;
        RECT 189.590 -41.090 190.040 -41.000 ;
        RECT 190.420 -41.100 190.870 -41.000 ;
        RECT 202.260 -40.750 202.710 -40.740 ;
        RECT 203.090 -40.750 203.540 -40.660 ;
        RECT 203.920 -40.740 205.450 -40.530 ;
        RECT 214.680 -40.530 215.130 -40.250 ;
        RECT 214.680 -40.740 216.210 -40.530 ;
        RECT 203.920 -40.750 204.370 -40.740 ;
        RECT 202.260 -41.000 204.370 -40.750 ;
        RECT 202.260 -41.100 202.710 -41.000 ;
        RECT 203.090 -41.090 203.540 -41.000 ;
        RECT 203.920 -41.100 204.370 -41.000 ;
        RECT 215.760 -40.750 216.210 -40.740 ;
        RECT 216.590 -40.730 217.030 -40.660 ;
        RECT 216.590 -40.750 217.690 -40.730 ;
        RECT 215.760 -41.000 217.690 -40.750 ;
        RECT 215.760 -41.100 216.210 -41.000 ;
        RECT 216.590 -41.050 217.690 -41.000 ;
        RECT 216.590 -41.090 217.030 -41.050 ;
      LAYER mcon ;
        RECT 12.270 16.370 12.530 16.630 ;
        RECT 16.100 16.370 16.360 16.630 ;
        RECT 25.770 16.370 26.030 16.630 ;
        RECT 29.600 16.370 29.860 16.630 ;
        RECT 39.270 16.370 39.530 16.630 ;
        RECT 43.100 16.370 43.360 16.630 ;
        RECT 52.770 16.370 53.030 16.630 ;
        RECT 56.600 16.370 56.860 16.630 ;
        RECT 12.270 13.540 12.530 13.800 ;
        RECT 16.100 13.540 16.360 13.800 ;
        RECT 66.270 16.370 66.530 16.630 ;
        RECT 70.100 16.370 70.360 16.630 ;
        RECT 25.770 13.540 26.030 13.800 ;
        RECT 29.600 13.540 29.860 13.800 ;
        RECT 79.770 16.370 80.030 16.630 ;
        RECT 83.600 16.370 83.860 16.630 ;
        RECT 39.270 13.540 39.530 13.800 ;
        RECT 43.100 13.540 43.360 13.800 ;
        RECT 93.270 16.370 93.530 16.630 ;
        RECT 97.100 16.370 97.360 16.630 ;
        RECT 52.770 13.540 53.030 13.800 ;
        RECT 56.600 13.540 56.860 13.800 ;
        RECT 106.770 16.370 107.030 16.630 ;
        RECT 110.600 16.370 110.860 16.630 ;
        RECT 66.270 13.540 66.530 13.800 ;
        RECT 70.100 13.540 70.360 13.800 ;
        RECT 120.270 16.370 120.530 16.630 ;
        RECT 124.100 16.370 124.360 16.630 ;
        RECT 79.770 13.540 80.030 13.800 ;
        RECT 83.600 13.540 83.860 13.800 ;
        RECT 133.770 16.370 134.030 16.630 ;
        RECT 137.600 16.370 137.860 16.630 ;
        RECT 93.270 13.540 93.530 13.800 ;
        RECT 97.100 13.540 97.360 13.800 ;
        RECT 147.270 16.370 147.530 16.630 ;
        RECT 151.100 16.370 151.360 16.630 ;
        RECT 106.770 13.540 107.030 13.800 ;
        RECT 110.600 13.540 110.860 13.800 ;
        RECT 160.770 16.370 161.030 16.630 ;
        RECT 164.600 16.370 164.860 16.630 ;
        RECT 120.270 13.540 120.530 13.800 ;
        RECT 124.100 13.540 124.360 13.800 ;
        RECT 174.270 16.370 174.530 16.630 ;
        RECT 178.100 16.370 178.360 16.630 ;
        RECT 133.770 13.540 134.030 13.800 ;
        RECT 137.600 13.540 137.860 13.800 ;
        RECT 187.770 16.370 188.030 16.630 ;
        RECT 191.600 16.370 191.860 16.630 ;
        RECT 147.270 13.540 147.530 13.800 ;
        RECT 151.100 13.540 151.360 13.800 ;
        RECT 201.270 16.370 201.530 16.630 ;
        RECT 205.100 16.370 205.360 16.630 ;
        RECT 160.770 13.540 161.030 13.800 ;
        RECT 164.600 13.540 164.860 13.800 ;
        RECT 214.770 16.370 215.030 16.630 ;
        RECT 174.270 13.540 174.530 13.800 ;
        RECT 178.100 13.540 178.360 13.800 ;
        RECT 187.770 13.540 188.030 13.800 ;
        RECT 191.600 13.540 191.860 13.800 ;
        RECT 201.270 13.540 201.530 13.800 ;
        RECT 205.100 13.540 205.360 13.800 ;
        RECT 214.770 13.540 215.030 13.800 ;
        RECT 12.270 12.760 12.530 13.020 ;
        RECT 16.100 12.760 16.360 13.020 ;
        RECT 25.770 12.760 26.030 13.020 ;
        RECT 29.600 12.760 29.860 13.020 ;
        RECT 39.270 12.760 39.530 13.020 ;
        RECT 43.100 12.760 43.360 13.020 ;
        RECT 52.770 12.760 53.030 13.020 ;
        RECT 56.600 12.760 56.860 13.020 ;
        RECT 12.270 9.930 12.530 10.190 ;
        RECT 16.100 9.930 16.360 10.190 ;
        RECT 66.270 12.760 66.530 13.020 ;
        RECT 70.100 12.760 70.360 13.020 ;
        RECT 25.770 9.930 26.030 10.190 ;
        RECT 29.600 9.930 29.860 10.190 ;
        RECT 79.770 12.760 80.030 13.020 ;
        RECT 83.600 12.760 83.860 13.020 ;
        RECT 39.270 9.930 39.530 10.190 ;
        RECT 43.100 9.930 43.360 10.190 ;
        RECT 93.270 12.760 93.530 13.020 ;
        RECT 97.100 12.760 97.360 13.020 ;
        RECT 52.770 9.930 53.030 10.190 ;
        RECT 56.600 9.930 56.860 10.190 ;
        RECT 106.770 12.760 107.030 13.020 ;
        RECT 110.600 12.760 110.860 13.020 ;
        RECT 66.270 9.930 66.530 10.190 ;
        RECT 70.100 9.930 70.360 10.190 ;
        RECT 120.270 12.760 120.530 13.020 ;
        RECT 124.100 12.760 124.360 13.020 ;
        RECT 79.770 9.930 80.030 10.190 ;
        RECT 83.600 9.930 83.860 10.190 ;
        RECT 133.770 12.760 134.030 13.020 ;
        RECT 137.600 12.760 137.860 13.020 ;
        RECT 93.270 9.930 93.530 10.190 ;
        RECT 97.100 9.930 97.360 10.190 ;
        RECT 147.270 12.760 147.530 13.020 ;
        RECT 151.100 12.760 151.360 13.020 ;
        RECT 106.770 9.930 107.030 10.190 ;
        RECT 110.600 9.930 110.860 10.190 ;
        RECT 160.770 12.760 161.030 13.020 ;
        RECT 164.600 12.760 164.860 13.020 ;
        RECT 120.270 9.930 120.530 10.190 ;
        RECT 124.100 9.930 124.360 10.190 ;
        RECT 174.270 12.760 174.530 13.020 ;
        RECT 178.100 12.760 178.360 13.020 ;
        RECT 133.770 9.930 134.030 10.190 ;
        RECT 137.600 9.930 137.860 10.190 ;
        RECT 187.770 12.760 188.030 13.020 ;
        RECT 191.600 12.760 191.860 13.020 ;
        RECT 147.270 9.930 147.530 10.190 ;
        RECT 151.100 9.930 151.360 10.190 ;
        RECT 201.270 12.760 201.530 13.020 ;
        RECT 205.100 12.760 205.360 13.020 ;
        RECT 160.770 9.930 161.030 10.190 ;
        RECT 164.600 9.930 164.860 10.190 ;
        RECT 214.770 12.760 215.030 13.020 ;
        RECT 174.270 9.930 174.530 10.190 ;
        RECT 178.100 9.930 178.360 10.190 ;
        RECT 187.770 9.930 188.030 10.190 ;
        RECT 191.600 9.930 191.860 10.190 ;
        RECT 201.270 9.930 201.530 10.190 ;
        RECT 205.100 9.930 205.360 10.190 ;
        RECT 214.770 9.930 215.030 10.190 ;
        RECT 12.270 9.150 12.530 9.410 ;
        RECT 16.100 9.150 16.360 9.410 ;
        RECT 25.770 9.150 26.030 9.410 ;
        RECT 29.600 9.150 29.860 9.410 ;
        RECT 39.270 9.150 39.530 9.410 ;
        RECT 43.100 9.150 43.360 9.410 ;
        RECT 52.770 9.150 53.030 9.410 ;
        RECT 56.600 9.150 56.860 9.410 ;
        RECT 12.270 6.320 12.530 6.580 ;
        RECT 16.100 6.320 16.360 6.580 ;
        RECT 66.270 9.150 66.530 9.410 ;
        RECT 70.100 9.150 70.360 9.410 ;
        RECT 25.770 6.320 26.030 6.580 ;
        RECT 29.600 6.320 29.860 6.580 ;
        RECT 79.770 9.150 80.030 9.410 ;
        RECT 83.600 9.150 83.860 9.410 ;
        RECT 39.270 6.320 39.530 6.580 ;
        RECT 43.100 6.320 43.360 6.580 ;
        RECT 93.270 9.150 93.530 9.410 ;
        RECT 97.100 9.150 97.360 9.410 ;
        RECT 52.770 6.320 53.030 6.580 ;
        RECT 56.600 6.320 56.860 6.580 ;
        RECT 106.770 9.150 107.030 9.410 ;
        RECT 110.600 9.150 110.860 9.410 ;
        RECT 66.270 6.320 66.530 6.580 ;
        RECT 70.100 6.320 70.360 6.580 ;
        RECT 120.270 9.150 120.530 9.410 ;
        RECT 124.100 9.150 124.360 9.410 ;
        RECT 79.770 6.320 80.030 6.580 ;
        RECT 83.600 6.320 83.860 6.580 ;
        RECT 133.770 9.150 134.030 9.410 ;
        RECT 137.600 9.150 137.860 9.410 ;
        RECT 93.270 6.320 93.530 6.580 ;
        RECT 97.100 6.320 97.360 6.580 ;
        RECT 147.270 9.150 147.530 9.410 ;
        RECT 151.100 9.150 151.360 9.410 ;
        RECT 106.770 6.320 107.030 6.580 ;
        RECT 110.600 6.320 110.860 6.580 ;
        RECT 160.770 9.150 161.030 9.410 ;
        RECT 164.600 9.150 164.860 9.410 ;
        RECT 120.270 6.320 120.530 6.580 ;
        RECT 124.100 6.320 124.360 6.580 ;
        RECT 174.270 9.150 174.530 9.410 ;
        RECT 178.100 9.150 178.360 9.410 ;
        RECT 133.770 6.320 134.030 6.580 ;
        RECT 137.600 6.320 137.860 6.580 ;
        RECT 187.770 9.150 188.030 9.410 ;
        RECT 191.600 9.150 191.860 9.410 ;
        RECT 147.270 6.320 147.530 6.580 ;
        RECT 151.100 6.320 151.360 6.580 ;
        RECT 201.270 9.150 201.530 9.410 ;
        RECT 205.100 9.150 205.360 9.410 ;
        RECT 160.770 6.320 161.030 6.580 ;
        RECT 164.600 6.320 164.860 6.580 ;
        RECT 214.770 9.150 215.030 9.410 ;
        RECT 174.270 6.320 174.530 6.580 ;
        RECT 178.100 6.320 178.360 6.580 ;
        RECT 187.770 6.320 188.030 6.580 ;
        RECT 191.600 6.320 191.860 6.580 ;
        RECT 201.270 6.320 201.530 6.580 ;
        RECT 205.100 6.320 205.360 6.580 ;
        RECT 214.770 6.320 215.030 6.580 ;
        RECT 12.270 5.540 12.530 5.800 ;
        RECT 16.100 5.540 16.360 5.800 ;
        RECT 25.770 5.540 26.030 5.800 ;
        RECT 29.600 5.540 29.860 5.800 ;
        RECT 39.270 5.540 39.530 5.800 ;
        RECT 43.100 5.540 43.360 5.800 ;
        RECT 52.770 5.540 53.030 5.800 ;
        RECT 56.600 5.540 56.860 5.800 ;
        RECT 12.270 2.710 12.530 2.970 ;
        RECT 16.100 2.710 16.360 2.970 ;
        RECT 66.270 5.540 66.530 5.800 ;
        RECT 70.100 5.540 70.360 5.800 ;
        RECT 25.770 2.710 26.030 2.970 ;
        RECT 29.600 2.710 29.860 2.970 ;
        RECT 79.770 5.540 80.030 5.800 ;
        RECT 83.600 5.540 83.860 5.800 ;
        RECT 39.270 2.710 39.530 2.970 ;
        RECT 43.100 2.710 43.360 2.970 ;
        RECT 93.270 5.540 93.530 5.800 ;
        RECT 97.100 5.540 97.360 5.800 ;
        RECT 52.770 2.710 53.030 2.970 ;
        RECT 56.600 2.710 56.860 2.970 ;
        RECT 106.770 5.540 107.030 5.800 ;
        RECT 110.600 5.540 110.860 5.800 ;
        RECT 66.270 2.710 66.530 2.970 ;
        RECT 70.100 2.710 70.360 2.970 ;
        RECT 120.270 5.540 120.530 5.800 ;
        RECT 124.100 5.540 124.360 5.800 ;
        RECT 79.770 2.710 80.030 2.970 ;
        RECT 83.600 2.710 83.860 2.970 ;
        RECT 133.770 5.540 134.030 5.800 ;
        RECT 137.600 5.540 137.860 5.800 ;
        RECT 93.270 2.710 93.530 2.970 ;
        RECT 97.100 2.710 97.360 2.970 ;
        RECT 147.270 5.540 147.530 5.800 ;
        RECT 151.100 5.540 151.360 5.800 ;
        RECT 106.770 2.710 107.030 2.970 ;
        RECT 110.600 2.710 110.860 2.970 ;
        RECT 160.770 5.540 161.030 5.800 ;
        RECT 164.600 5.540 164.860 5.800 ;
        RECT 120.270 2.710 120.530 2.970 ;
        RECT 124.100 2.710 124.360 2.970 ;
        RECT 174.270 5.540 174.530 5.800 ;
        RECT 178.100 5.540 178.360 5.800 ;
        RECT 133.770 2.710 134.030 2.970 ;
        RECT 137.600 2.710 137.860 2.970 ;
        RECT 187.770 5.540 188.030 5.800 ;
        RECT 191.600 5.540 191.860 5.800 ;
        RECT 147.270 2.710 147.530 2.970 ;
        RECT 151.100 2.710 151.360 2.970 ;
        RECT 201.270 5.540 201.530 5.800 ;
        RECT 205.100 5.540 205.360 5.800 ;
        RECT 160.770 2.710 161.030 2.970 ;
        RECT 164.600 2.710 164.860 2.970 ;
        RECT 214.770 5.540 215.030 5.800 ;
        RECT 174.270 2.710 174.530 2.970 ;
        RECT 178.100 2.710 178.360 2.970 ;
        RECT 187.770 2.710 188.030 2.970 ;
        RECT 191.600 2.710 191.860 2.970 ;
        RECT 201.270 2.710 201.530 2.970 ;
        RECT 205.100 2.710 205.360 2.970 ;
        RECT 214.770 2.710 215.030 2.970 ;
        RECT 12.270 1.930 12.530 2.190 ;
        RECT 16.100 1.930 16.360 2.190 ;
        RECT 25.770 1.930 26.030 2.190 ;
        RECT 29.600 1.930 29.860 2.190 ;
        RECT 39.270 1.930 39.530 2.190 ;
        RECT 43.100 1.930 43.360 2.190 ;
        RECT 52.770 1.930 53.030 2.190 ;
        RECT 56.600 1.930 56.860 2.190 ;
        RECT 12.270 -0.900 12.530 -0.640 ;
        RECT 16.100 -0.900 16.360 -0.640 ;
        RECT 66.270 1.930 66.530 2.190 ;
        RECT 70.100 1.930 70.360 2.190 ;
        RECT 25.770 -0.900 26.030 -0.640 ;
        RECT 29.600 -0.900 29.860 -0.640 ;
        RECT 79.770 1.930 80.030 2.190 ;
        RECT 83.600 1.930 83.860 2.190 ;
        RECT 39.270 -0.900 39.530 -0.640 ;
        RECT 43.100 -0.900 43.360 -0.640 ;
        RECT 93.270 1.930 93.530 2.190 ;
        RECT 97.100 1.930 97.360 2.190 ;
        RECT 52.770 -0.900 53.030 -0.640 ;
        RECT 56.600 -0.900 56.860 -0.640 ;
        RECT 106.770 1.930 107.030 2.190 ;
        RECT 110.600 1.930 110.860 2.190 ;
        RECT 66.270 -0.900 66.530 -0.640 ;
        RECT 70.100 -0.900 70.360 -0.640 ;
        RECT 120.270 1.930 120.530 2.190 ;
        RECT 124.100 1.930 124.360 2.190 ;
        RECT 79.770 -0.900 80.030 -0.640 ;
        RECT 83.600 -0.900 83.860 -0.640 ;
        RECT 133.770 1.930 134.030 2.190 ;
        RECT 137.600 1.930 137.860 2.190 ;
        RECT 93.270 -0.900 93.530 -0.640 ;
        RECT 97.100 -0.900 97.360 -0.640 ;
        RECT 147.270 1.930 147.530 2.190 ;
        RECT 151.100 1.930 151.360 2.190 ;
        RECT 106.770 -0.900 107.030 -0.640 ;
        RECT 110.600 -0.900 110.860 -0.640 ;
        RECT 160.770 1.930 161.030 2.190 ;
        RECT 164.600 1.930 164.860 2.190 ;
        RECT 120.270 -0.900 120.530 -0.640 ;
        RECT 124.100 -0.900 124.360 -0.640 ;
        RECT 174.270 1.930 174.530 2.190 ;
        RECT 178.100 1.930 178.360 2.190 ;
        RECT 133.770 -0.900 134.030 -0.640 ;
        RECT 137.600 -0.900 137.860 -0.640 ;
        RECT 187.770 1.930 188.030 2.190 ;
        RECT 191.600 1.930 191.860 2.190 ;
        RECT 147.270 -0.900 147.530 -0.640 ;
        RECT 151.100 -0.900 151.360 -0.640 ;
        RECT 201.270 1.930 201.530 2.190 ;
        RECT 205.100 1.930 205.360 2.190 ;
        RECT 160.770 -0.900 161.030 -0.640 ;
        RECT 164.600 -0.900 164.860 -0.640 ;
        RECT 214.770 1.930 215.030 2.190 ;
        RECT 174.270 -0.900 174.530 -0.640 ;
        RECT 178.100 -0.900 178.360 -0.640 ;
        RECT 187.770 -0.900 188.030 -0.640 ;
        RECT 191.600 -0.900 191.860 -0.640 ;
        RECT 201.270 -0.900 201.530 -0.640 ;
        RECT 205.100 -0.900 205.360 -0.640 ;
        RECT 214.770 -0.900 215.030 -0.640 ;
        RECT 12.270 -1.680 12.530 -1.420 ;
        RECT 16.100 -1.680 16.360 -1.420 ;
        RECT 25.770 -1.680 26.030 -1.420 ;
        RECT 29.600 -1.680 29.860 -1.420 ;
        RECT 39.270 -1.680 39.530 -1.420 ;
        RECT 43.100 -1.680 43.360 -1.420 ;
        RECT 52.770 -1.680 53.030 -1.420 ;
        RECT 56.600 -1.680 56.860 -1.420 ;
        RECT 12.270 -4.510 12.530 -4.250 ;
        RECT 16.100 -4.510 16.360 -4.250 ;
        RECT 66.270 -1.680 66.530 -1.420 ;
        RECT 70.100 -1.680 70.360 -1.420 ;
        RECT 25.770 -4.510 26.030 -4.250 ;
        RECT 29.600 -4.510 29.860 -4.250 ;
        RECT 79.770 -1.680 80.030 -1.420 ;
        RECT 83.600 -1.680 83.860 -1.420 ;
        RECT 39.270 -4.510 39.530 -4.250 ;
        RECT 43.100 -4.510 43.360 -4.250 ;
        RECT 93.270 -1.680 93.530 -1.420 ;
        RECT 97.100 -1.680 97.360 -1.420 ;
        RECT 52.770 -4.510 53.030 -4.250 ;
        RECT 56.600 -4.510 56.860 -4.250 ;
        RECT 106.770 -1.680 107.030 -1.420 ;
        RECT 110.600 -1.680 110.860 -1.420 ;
        RECT 66.270 -4.510 66.530 -4.250 ;
        RECT 70.100 -4.510 70.360 -4.250 ;
        RECT 120.270 -1.680 120.530 -1.420 ;
        RECT 124.100 -1.680 124.360 -1.420 ;
        RECT 79.770 -4.510 80.030 -4.250 ;
        RECT 83.600 -4.510 83.860 -4.250 ;
        RECT 133.770 -1.680 134.030 -1.420 ;
        RECT 137.600 -1.680 137.860 -1.420 ;
        RECT 93.270 -4.510 93.530 -4.250 ;
        RECT 97.100 -4.510 97.360 -4.250 ;
        RECT 147.270 -1.680 147.530 -1.420 ;
        RECT 151.100 -1.680 151.360 -1.420 ;
        RECT 106.770 -4.510 107.030 -4.250 ;
        RECT 110.600 -4.510 110.860 -4.250 ;
        RECT 160.770 -1.680 161.030 -1.420 ;
        RECT 164.600 -1.680 164.860 -1.420 ;
        RECT 120.270 -4.510 120.530 -4.250 ;
        RECT 124.100 -4.510 124.360 -4.250 ;
        RECT 174.270 -1.680 174.530 -1.420 ;
        RECT 178.100 -1.680 178.360 -1.420 ;
        RECT 133.770 -4.510 134.030 -4.250 ;
        RECT 137.600 -4.510 137.860 -4.250 ;
        RECT 187.770 -1.680 188.030 -1.420 ;
        RECT 191.600 -1.680 191.860 -1.420 ;
        RECT 147.270 -4.510 147.530 -4.250 ;
        RECT 151.100 -4.510 151.360 -4.250 ;
        RECT 201.270 -1.680 201.530 -1.420 ;
        RECT 205.100 -1.680 205.360 -1.420 ;
        RECT 160.770 -4.510 161.030 -4.250 ;
        RECT 164.600 -4.510 164.860 -4.250 ;
        RECT 214.770 -1.680 215.030 -1.420 ;
        RECT 174.270 -4.510 174.530 -4.250 ;
        RECT 178.100 -4.510 178.360 -4.250 ;
        RECT 187.770 -4.510 188.030 -4.250 ;
        RECT 191.600 -4.510 191.860 -4.250 ;
        RECT 201.270 -4.510 201.530 -4.250 ;
        RECT 205.100 -4.510 205.360 -4.250 ;
        RECT 214.770 -4.510 215.030 -4.250 ;
        RECT 12.270 -5.290 12.530 -5.030 ;
        RECT 16.100 -5.290 16.360 -5.030 ;
        RECT 25.770 -5.290 26.030 -5.030 ;
        RECT 29.600 -5.290 29.860 -5.030 ;
        RECT 39.270 -5.290 39.530 -5.030 ;
        RECT 43.100 -5.290 43.360 -5.030 ;
        RECT 52.770 -5.290 53.030 -5.030 ;
        RECT 56.600 -5.290 56.860 -5.030 ;
        RECT 12.270 -8.120 12.530 -7.860 ;
        RECT 16.100 -8.120 16.360 -7.860 ;
        RECT 66.270 -5.290 66.530 -5.030 ;
        RECT 70.100 -5.290 70.360 -5.030 ;
        RECT 25.770 -8.120 26.030 -7.860 ;
        RECT 29.600 -8.120 29.860 -7.860 ;
        RECT 79.770 -5.290 80.030 -5.030 ;
        RECT 83.600 -5.290 83.860 -5.030 ;
        RECT 39.270 -8.120 39.530 -7.860 ;
        RECT 43.100 -8.120 43.360 -7.860 ;
        RECT 93.270 -5.290 93.530 -5.030 ;
        RECT 97.100 -5.290 97.360 -5.030 ;
        RECT 52.770 -8.120 53.030 -7.860 ;
        RECT 56.600 -8.120 56.860 -7.860 ;
        RECT 106.770 -5.290 107.030 -5.030 ;
        RECT 110.600 -5.290 110.860 -5.030 ;
        RECT 66.270 -8.120 66.530 -7.860 ;
        RECT 70.100 -8.120 70.360 -7.860 ;
        RECT 120.270 -5.290 120.530 -5.030 ;
        RECT 124.100 -5.290 124.360 -5.030 ;
        RECT 79.770 -8.120 80.030 -7.860 ;
        RECT 83.600 -8.120 83.860 -7.860 ;
        RECT 133.770 -5.290 134.030 -5.030 ;
        RECT 137.600 -5.290 137.860 -5.030 ;
        RECT 93.270 -8.120 93.530 -7.860 ;
        RECT 97.100 -8.120 97.360 -7.860 ;
        RECT 147.270 -5.290 147.530 -5.030 ;
        RECT 151.100 -5.290 151.360 -5.030 ;
        RECT 106.770 -8.120 107.030 -7.860 ;
        RECT 110.600 -8.120 110.860 -7.860 ;
        RECT 160.770 -5.290 161.030 -5.030 ;
        RECT 164.600 -5.290 164.860 -5.030 ;
        RECT 120.270 -8.120 120.530 -7.860 ;
        RECT 124.100 -8.120 124.360 -7.860 ;
        RECT 174.270 -5.290 174.530 -5.030 ;
        RECT 178.100 -5.290 178.360 -5.030 ;
        RECT 133.770 -8.120 134.030 -7.860 ;
        RECT 137.600 -8.120 137.860 -7.860 ;
        RECT 187.770 -5.290 188.030 -5.030 ;
        RECT 191.600 -5.290 191.860 -5.030 ;
        RECT 147.270 -8.120 147.530 -7.860 ;
        RECT 151.100 -8.120 151.360 -7.860 ;
        RECT 201.270 -5.290 201.530 -5.030 ;
        RECT 205.100 -5.290 205.360 -5.030 ;
        RECT 160.770 -8.120 161.030 -7.860 ;
        RECT 164.600 -8.120 164.860 -7.860 ;
        RECT 214.770 -5.290 215.030 -5.030 ;
        RECT 174.270 -8.120 174.530 -7.860 ;
        RECT 178.100 -8.120 178.360 -7.860 ;
        RECT 187.770 -8.120 188.030 -7.860 ;
        RECT 191.600 -8.120 191.860 -7.860 ;
        RECT 201.270 -8.120 201.530 -7.860 ;
        RECT 205.100 -8.120 205.360 -7.860 ;
        RECT 214.770 -8.120 215.030 -7.860 ;
        RECT 12.270 -8.900 12.530 -8.640 ;
        RECT 16.100 -8.900 16.360 -8.640 ;
        RECT 25.770 -8.900 26.030 -8.640 ;
        RECT 29.600 -8.900 29.860 -8.640 ;
        RECT 39.270 -8.900 39.530 -8.640 ;
        RECT 43.100 -8.900 43.360 -8.640 ;
        RECT 52.770 -8.900 53.030 -8.640 ;
        RECT 56.600 -8.900 56.860 -8.640 ;
        RECT 12.270 -11.730 12.530 -11.470 ;
        RECT 16.100 -11.730 16.360 -11.470 ;
        RECT 66.270 -8.900 66.530 -8.640 ;
        RECT 70.100 -8.900 70.360 -8.640 ;
        RECT 25.770 -11.730 26.030 -11.470 ;
        RECT 29.600 -11.730 29.860 -11.470 ;
        RECT 79.770 -8.900 80.030 -8.640 ;
        RECT 83.600 -8.900 83.860 -8.640 ;
        RECT 39.270 -11.730 39.530 -11.470 ;
        RECT 43.100 -11.730 43.360 -11.470 ;
        RECT 93.270 -8.900 93.530 -8.640 ;
        RECT 97.100 -8.900 97.360 -8.640 ;
        RECT 52.770 -11.730 53.030 -11.470 ;
        RECT 56.600 -11.730 56.860 -11.470 ;
        RECT 106.770 -8.900 107.030 -8.640 ;
        RECT 110.600 -8.900 110.860 -8.640 ;
        RECT 66.270 -11.730 66.530 -11.470 ;
        RECT 70.100 -11.730 70.360 -11.470 ;
        RECT 120.270 -8.900 120.530 -8.640 ;
        RECT 124.100 -8.900 124.360 -8.640 ;
        RECT 79.770 -11.730 80.030 -11.470 ;
        RECT 83.600 -11.730 83.860 -11.470 ;
        RECT 133.770 -8.900 134.030 -8.640 ;
        RECT 137.600 -8.900 137.860 -8.640 ;
        RECT 93.270 -11.730 93.530 -11.470 ;
        RECT 97.100 -11.730 97.360 -11.470 ;
        RECT 147.270 -8.900 147.530 -8.640 ;
        RECT 151.100 -8.900 151.360 -8.640 ;
        RECT 106.770 -11.730 107.030 -11.470 ;
        RECT 110.600 -11.730 110.860 -11.470 ;
        RECT 160.770 -8.900 161.030 -8.640 ;
        RECT 164.600 -8.900 164.860 -8.640 ;
        RECT 120.270 -11.730 120.530 -11.470 ;
        RECT 124.100 -11.730 124.360 -11.470 ;
        RECT 174.270 -8.900 174.530 -8.640 ;
        RECT 178.100 -8.900 178.360 -8.640 ;
        RECT 133.770 -11.730 134.030 -11.470 ;
        RECT 137.600 -11.730 137.860 -11.470 ;
        RECT 187.770 -8.900 188.030 -8.640 ;
        RECT 191.600 -8.900 191.860 -8.640 ;
        RECT 147.270 -11.730 147.530 -11.470 ;
        RECT 151.100 -11.730 151.360 -11.470 ;
        RECT 201.270 -8.900 201.530 -8.640 ;
        RECT 205.100 -8.900 205.360 -8.640 ;
        RECT 160.770 -11.730 161.030 -11.470 ;
        RECT 164.600 -11.730 164.860 -11.470 ;
        RECT 214.770 -8.900 215.030 -8.640 ;
        RECT 174.270 -11.730 174.530 -11.470 ;
        RECT 178.100 -11.730 178.360 -11.470 ;
        RECT 187.770 -11.730 188.030 -11.470 ;
        RECT 191.600 -11.730 191.860 -11.470 ;
        RECT 201.270 -11.730 201.530 -11.470 ;
        RECT 205.100 -11.730 205.360 -11.470 ;
        RECT 214.770 -11.730 215.030 -11.470 ;
        RECT 12.270 -12.510 12.530 -12.250 ;
        RECT 16.100 -12.510 16.360 -12.250 ;
        RECT 25.770 -12.510 26.030 -12.250 ;
        RECT 29.600 -12.510 29.860 -12.250 ;
        RECT 39.270 -12.510 39.530 -12.250 ;
        RECT 43.100 -12.510 43.360 -12.250 ;
        RECT 52.770 -12.510 53.030 -12.250 ;
        RECT 56.600 -12.510 56.860 -12.250 ;
        RECT 12.270 -15.340 12.530 -15.080 ;
        RECT 16.100 -15.340 16.360 -15.080 ;
        RECT 66.270 -12.510 66.530 -12.250 ;
        RECT 70.100 -12.510 70.360 -12.250 ;
        RECT 25.770 -15.340 26.030 -15.080 ;
        RECT 29.600 -15.340 29.860 -15.080 ;
        RECT 79.770 -12.510 80.030 -12.250 ;
        RECT 83.600 -12.510 83.860 -12.250 ;
        RECT 39.270 -15.340 39.530 -15.080 ;
        RECT 43.100 -15.340 43.360 -15.080 ;
        RECT 93.270 -12.510 93.530 -12.250 ;
        RECT 97.100 -12.510 97.360 -12.250 ;
        RECT 52.770 -15.340 53.030 -15.080 ;
        RECT 56.600 -15.340 56.860 -15.080 ;
        RECT 106.770 -12.510 107.030 -12.250 ;
        RECT 110.600 -12.510 110.860 -12.250 ;
        RECT 66.270 -15.340 66.530 -15.080 ;
        RECT 70.100 -15.340 70.360 -15.080 ;
        RECT 120.270 -12.510 120.530 -12.250 ;
        RECT 124.100 -12.510 124.360 -12.250 ;
        RECT 79.770 -15.340 80.030 -15.080 ;
        RECT 83.600 -15.340 83.860 -15.080 ;
        RECT 133.770 -12.510 134.030 -12.250 ;
        RECT 137.600 -12.510 137.860 -12.250 ;
        RECT 93.270 -15.340 93.530 -15.080 ;
        RECT 97.100 -15.340 97.360 -15.080 ;
        RECT 147.270 -12.510 147.530 -12.250 ;
        RECT 151.100 -12.510 151.360 -12.250 ;
        RECT 106.770 -15.340 107.030 -15.080 ;
        RECT 110.600 -15.340 110.860 -15.080 ;
        RECT 160.770 -12.510 161.030 -12.250 ;
        RECT 164.600 -12.510 164.860 -12.250 ;
        RECT 120.270 -15.340 120.530 -15.080 ;
        RECT 124.100 -15.340 124.360 -15.080 ;
        RECT 174.270 -12.510 174.530 -12.250 ;
        RECT 178.100 -12.510 178.360 -12.250 ;
        RECT 133.770 -15.340 134.030 -15.080 ;
        RECT 137.600 -15.340 137.860 -15.080 ;
        RECT 187.770 -12.510 188.030 -12.250 ;
        RECT 191.600 -12.510 191.860 -12.250 ;
        RECT 147.270 -15.340 147.530 -15.080 ;
        RECT 151.100 -15.340 151.360 -15.080 ;
        RECT 201.270 -12.510 201.530 -12.250 ;
        RECT 205.100 -12.510 205.360 -12.250 ;
        RECT 160.770 -15.340 161.030 -15.080 ;
        RECT 164.600 -15.340 164.860 -15.080 ;
        RECT 214.770 -12.510 215.030 -12.250 ;
        RECT 174.270 -15.340 174.530 -15.080 ;
        RECT 178.100 -15.340 178.360 -15.080 ;
        RECT 187.770 -15.340 188.030 -15.080 ;
        RECT 191.600 -15.340 191.860 -15.080 ;
        RECT 201.270 -15.340 201.530 -15.080 ;
        RECT 205.100 -15.340 205.360 -15.080 ;
        RECT 214.770 -15.340 215.030 -15.080 ;
        RECT 12.270 -16.120 12.530 -15.860 ;
        RECT 16.100 -16.120 16.360 -15.860 ;
        RECT 25.770 -16.120 26.030 -15.860 ;
        RECT 29.600 -16.120 29.860 -15.860 ;
        RECT 39.270 -16.120 39.530 -15.860 ;
        RECT 43.100 -16.120 43.360 -15.860 ;
        RECT 52.770 -16.120 53.030 -15.860 ;
        RECT 56.600 -16.120 56.860 -15.860 ;
        RECT 12.270 -18.950 12.530 -18.690 ;
        RECT 16.100 -18.950 16.360 -18.690 ;
        RECT 66.270 -16.120 66.530 -15.860 ;
        RECT 70.100 -16.120 70.360 -15.860 ;
        RECT 25.770 -18.950 26.030 -18.690 ;
        RECT 29.600 -18.950 29.860 -18.690 ;
        RECT 79.770 -16.120 80.030 -15.860 ;
        RECT 83.600 -16.120 83.860 -15.860 ;
        RECT 39.270 -18.950 39.530 -18.690 ;
        RECT 43.100 -18.950 43.360 -18.690 ;
        RECT 93.270 -16.120 93.530 -15.860 ;
        RECT 97.100 -16.120 97.360 -15.860 ;
        RECT 52.770 -18.950 53.030 -18.690 ;
        RECT 56.600 -18.950 56.860 -18.690 ;
        RECT 106.770 -16.120 107.030 -15.860 ;
        RECT 110.600 -16.120 110.860 -15.860 ;
        RECT 66.270 -18.950 66.530 -18.690 ;
        RECT 70.100 -18.950 70.360 -18.690 ;
        RECT 120.270 -16.120 120.530 -15.860 ;
        RECT 124.100 -16.120 124.360 -15.860 ;
        RECT 79.770 -18.950 80.030 -18.690 ;
        RECT 83.600 -18.950 83.860 -18.690 ;
        RECT 133.770 -16.120 134.030 -15.860 ;
        RECT 137.600 -16.120 137.860 -15.860 ;
        RECT 93.270 -18.950 93.530 -18.690 ;
        RECT 97.100 -18.950 97.360 -18.690 ;
        RECT 147.270 -16.120 147.530 -15.860 ;
        RECT 151.100 -16.120 151.360 -15.860 ;
        RECT 106.770 -18.950 107.030 -18.690 ;
        RECT 110.600 -18.950 110.860 -18.690 ;
        RECT 160.770 -16.120 161.030 -15.860 ;
        RECT 164.600 -16.120 164.860 -15.860 ;
        RECT 120.270 -18.950 120.530 -18.690 ;
        RECT 124.100 -18.950 124.360 -18.690 ;
        RECT 174.270 -16.120 174.530 -15.860 ;
        RECT 178.100 -16.120 178.360 -15.860 ;
        RECT 133.770 -18.950 134.030 -18.690 ;
        RECT 137.600 -18.950 137.860 -18.690 ;
        RECT 187.770 -16.120 188.030 -15.860 ;
        RECT 191.600 -16.120 191.860 -15.860 ;
        RECT 147.270 -18.950 147.530 -18.690 ;
        RECT 151.100 -18.950 151.360 -18.690 ;
        RECT 201.270 -16.120 201.530 -15.860 ;
        RECT 205.100 -16.120 205.360 -15.860 ;
        RECT 160.770 -18.950 161.030 -18.690 ;
        RECT 164.600 -18.950 164.860 -18.690 ;
        RECT 214.770 -16.120 215.030 -15.860 ;
        RECT 174.270 -18.950 174.530 -18.690 ;
        RECT 178.100 -18.950 178.360 -18.690 ;
        RECT 187.770 -18.950 188.030 -18.690 ;
        RECT 191.600 -18.950 191.860 -18.690 ;
        RECT 201.270 -18.950 201.530 -18.690 ;
        RECT 205.100 -18.950 205.360 -18.690 ;
        RECT 214.770 -18.950 215.030 -18.690 ;
        RECT 12.270 -19.730 12.530 -19.470 ;
        RECT 16.100 -19.730 16.360 -19.470 ;
        RECT 25.770 -19.730 26.030 -19.470 ;
        RECT 29.600 -19.730 29.860 -19.470 ;
        RECT 39.270 -19.730 39.530 -19.470 ;
        RECT 43.100 -19.730 43.360 -19.470 ;
        RECT 52.770 -19.730 53.030 -19.470 ;
        RECT 56.600 -19.730 56.860 -19.470 ;
        RECT 12.270 -22.560 12.530 -22.300 ;
        RECT 16.100 -22.560 16.360 -22.300 ;
        RECT 66.270 -19.730 66.530 -19.470 ;
        RECT 70.100 -19.730 70.360 -19.470 ;
        RECT 25.770 -22.560 26.030 -22.300 ;
        RECT 29.600 -22.560 29.860 -22.300 ;
        RECT 79.770 -19.730 80.030 -19.470 ;
        RECT 83.600 -19.730 83.860 -19.470 ;
        RECT 39.270 -22.560 39.530 -22.300 ;
        RECT 43.100 -22.560 43.360 -22.300 ;
        RECT 93.270 -19.730 93.530 -19.470 ;
        RECT 97.100 -19.730 97.360 -19.470 ;
        RECT 52.770 -22.560 53.030 -22.300 ;
        RECT 56.600 -22.560 56.860 -22.300 ;
        RECT 106.770 -19.730 107.030 -19.470 ;
        RECT 110.600 -19.730 110.860 -19.470 ;
        RECT 66.270 -22.560 66.530 -22.300 ;
        RECT 70.100 -22.560 70.360 -22.300 ;
        RECT 120.270 -19.730 120.530 -19.470 ;
        RECT 124.100 -19.730 124.360 -19.470 ;
        RECT 79.770 -22.560 80.030 -22.300 ;
        RECT 83.600 -22.560 83.860 -22.300 ;
        RECT 133.770 -19.730 134.030 -19.470 ;
        RECT 137.600 -19.730 137.860 -19.470 ;
        RECT 93.270 -22.560 93.530 -22.300 ;
        RECT 97.100 -22.560 97.360 -22.300 ;
        RECT 147.270 -19.730 147.530 -19.470 ;
        RECT 151.100 -19.730 151.360 -19.470 ;
        RECT 106.770 -22.560 107.030 -22.300 ;
        RECT 110.600 -22.560 110.860 -22.300 ;
        RECT 160.770 -19.730 161.030 -19.470 ;
        RECT 164.600 -19.730 164.860 -19.470 ;
        RECT 120.270 -22.560 120.530 -22.300 ;
        RECT 124.100 -22.560 124.360 -22.300 ;
        RECT 174.270 -19.730 174.530 -19.470 ;
        RECT 178.100 -19.730 178.360 -19.470 ;
        RECT 133.770 -22.560 134.030 -22.300 ;
        RECT 137.600 -22.560 137.860 -22.300 ;
        RECT 187.770 -19.730 188.030 -19.470 ;
        RECT 191.600 -19.730 191.860 -19.470 ;
        RECT 147.270 -22.560 147.530 -22.300 ;
        RECT 151.100 -22.560 151.360 -22.300 ;
        RECT 201.270 -19.730 201.530 -19.470 ;
        RECT 205.100 -19.730 205.360 -19.470 ;
        RECT 160.770 -22.560 161.030 -22.300 ;
        RECT 164.600 -22.560 164.860 -22.300 ;
        RECT 214.770 -19.730 215.030 -19.470 ;
        RECT 174.270 -22.560 174.530 -22.300 ;
        RECT 178.100 -22.560 178.360 -22.300 ;
        RECT 187.770 -22.560 188.030 -22.300 ;
        RECT 191.600 -22.560 191.860 -22.300 ;
        RECT 201.270 -22.560 201.530 -22.300 ;
        RECT 205.100 -22.560 205.360 -22.300 ;
        RECT 214.770 -22.560 215.030 -22.300 ;
        RECT 12.270 -23.340 12.530 -23.080 ;
        RECT 16.100 -23.340 16.360 -23.080 ;
        RECT 25.770 -23.340 26.030 -23.080 ;
        RECT 29.600 -23.340 29.860 -23.080 ;
        RECT 39.270 -23.340 39.530 -23.080 ;
        RECT 43.100 -23.340 43.360 -23.080 ;
        RECT 52.770 -23.340 53.030 -23.080 ;
        RECT 56.600 -23.340 56.860 -23.080 ;
        RECT 12.270 -26.170 12.530 -25.910 ;
        RECT 16.100 -26.170 16.360 -25.910 ;
        RECT 66.270 -23.340 66.530 -23.080 ;
        RECT 70.100 -23.340 70.360 -23.080 ;
        RECT 25.770 -26.170 26.030 -25.910 ;
        RECT 29.600 -26.170 29.860 -25.910 ;
        RECT 79.770 -23.340 80.030 -23.080 ;
        RECT 83.600 -23.340 83.860 -23.080 ;
        RECT 39.270 -26.170 39.530 -25.910 ;
        RECT 43.100 -26.170 43.360 -25.910 ;
        RECT 93.270 -23.340 93.530 -23.080 ;
        RECT 97.100 -23.340 97.360 -23.080 ;
        RECT 52.770 -26.170 53.030 -25.910 ;
        RECT 56.600 -26.170 56.860 -25.910 ;
        RECT 106.770 -23.340 107.030 -23.080 ;
        RECT 110.600 -23.340 110.860 -23.080 ;
        RECT 66.270 -26.170 66.530 -25.910 ;
        RECT 70.100 -26.170 70.360 -25.910 ;
        RECT 120.270 -23.340 120.530 -23.080 ;
        RECT 124.100 -23.340 124.360 -23.080 ;
        RECT 79.770 -26.170 80.030 -25.910 ;
        RECT 83.600 -26.170 83.860 -25.910 ;
        RECT 133.770 -23.340 134.030 -23.080 ;
        RECT 137.600 -23.340 137.860 -23.080 ;
        RECT 93.270 -26.170 93.530 -25.910 ;
        RECT 97.100 -26.170 97.360 -25.910 ;
        RECT 147.270 -23.340 147.530 -23.080 ;
        RECT 151.100 -23.340 151.360 -23.080 ;
        RECT 106.770 -26.170 107.030 -25.910 ;
        RECT 110.600 -26.170 110.860 -25.910 ;
        RECT 160.770 -23.340 161.030 -23.080 ;
        RECT 164.600 -23.340 164.860 -23.080 ;
        RECT 120.270 -26.170 120.530 -25.910 ;
        RECT 124.100 -26.170 124.360 -25.910 ;
        RECT 174.270 -23.340 174.530 -23.080 ;
        RECT 178.100 -23.340 178.360 -23.080 ;
        RECT 133.770 -26.170 134.030 -25.910 ;
        RECT 137.600 -26.170 137.860 -25.910 ;
        RECT 187.770 -23.340 188.030 -23.080 ;
        RECT 191.600 -23.340 191.860 -23.080 ;
        RECT 147.270 -26.170 147.530 -25.910 ;
        RECT 151.100 -26.170 151.360 -25.910 ;
        RECT 201.270 -23.340 201.530 -23.080 ;
        RECT 205.100 -23.340 205.360 -23.080 ;
        RECT 160.770 -26.170 161.030 -25.910 ;
        RECT 164.600 -26.170 164.860 -25.910 ;
        RECT 214.770 -23.340 215.030 -23.080 ;
        RECT 174.270 -26.170 174.530 -25.910 ;
        RECT 178.100 -26.170 178.360 -25.910 ;
        RECT 187.770 -26.170 188.030 -25.910 ;
        RECT 191.600 -26.170 191.860 -25.910 ;
        RECT 201.270 -26.170 201.530 -25.910 ;
        RECT 205.100 -26.170 205.360 -25.910 ;
        RECT 214.770 -26.170 215.030 -25.910 ;
        RECT 12.270 -26.950 12.530 -26.690 ;
        RECT 16.100 -26.950 16.360 -26.690 ;
        RECT 25.770 -26.950 26.030 -26.690 ;
        RECT 29.600 -26.950 29.860 -26.690 ;
        RECT 39.270 -26.950 39.530 -26.690 ;
        RECT 43.100 -26.950 43.360 -26.690 ;
        RECT 52.770 -26.950 53.030 -26.690 ;
        RECT 56.600 -26.950 56.860 -26.690 ;
        RECT 12.270 -29.780 12.530 -29.520 ;
        RECT 16.100 -29.780 16.360 -29.520 ;
        RECT 66.270 -26.950 66.530 -26.690 ;
        RECT 70.100 -26.950 70.360 -26.690 ;
        RECT 25.770 -29.780 26.030 -29.520 ;
        RECT 29.600 -29.780 29.860 -29.520 ;
        RECT 79.770 -26.950 80.030 -26.690 ;
        RECT 83.600 -26.950 83.860 -26.690 ;
        RECT 39.270 -29.780 39.530 -29.520 ;
        RECT 43.100 -29.780 43.360 -29.520 ;
        RECT 93.270 -26.950 93.530 -26.690 ;
        RECT 97.100 -26.950 97.360 -26.690 ;
        RECT 52.770 -29.780 53.030 -29.520 ;
        RECT 56.600 -29.780 56.860 -29.520 ;
        RECT 106.770 -26.950 107.030 -26.690 ;
        RECT 110.600 -26.950 110.860 -26.690 ;
        RECT 66.270 -29.780 66.530 -29.520 ;
        RECT 70.100 -29.780 70.360 -29.520 ;
        RECT 120.270 -26.950 120.530 -26.690 ;
        RECT 124.100 -26.950 124.360 -26.690 ;
        RECT 79.770 -29.780 80.030 -29.520 ;
        RECT 83.600 -29.780 83.860 -29.520 ;
        RECT 133.770 -26.950 134.030 -26.690 ;
        RECT 137.600 -26.950 137.860 -26.690 ;
        RECT 93.270 -29.780 93.530 -29.520 ;
        RECT 97.100 -29.780 97.360 -29.520 ;
        RECT 147.270 -26.950 147.530 -26.690 ;
        RECT 151.100 -26.950 151.360 -26.690 ;
        RECT 106.770 -29.780 107.030 -29.520 ;
        RECT 110.600 -29.780 110.860 -29.520 ;
        RECT 160.770 -26.950 161.030 -26.690 ;
        RECT 164.600 -26.950 164.860 -26.690 ;
        RECT 120.270 -29.780 120.530 -29.520 ;
        RECT 124.100 -29.780 124.360 -29.520 ;
        RECT 174.270 -26.950 174.530 -26.690 ;
        RECT 178.100 -26.950 178.360 -26.690 ;
        RECT 133.770 -29.780 134.030 -29.520 ;
        RECT 137.600 -29.780 137.860 -29.520 ;
        RECT 187.770 -26.950 188.030 -26.690 ;
        RECT 191.600 -26.950 191.860 -26.690 ;
        RECT 147.270 -29.780 147.530 -29.520 ;
        RECT 151.100 -29.780 151.360 -29.520 ;
        RECT 201.270 -26.950 201.530 -26.690 ;
        RECT 205.100 -26.950 205.360 -26.690 ;
        RECT 160.770 -29.780 161.030 -29.520 ;
        RECT 164.600 -29.780 164.860 -29.520 ;
        RECT 214.770 -26.950 215.030 -26.690 ;
        RECT 174.270 -29.780 174.530 -29.520 ;
        RECT 178.100 -29.780 178.360 -29.520 ;
        RECT 187.770 -29.780 188.030 -29.520 ;
        RECT 191.600 -29.780 191.860 -29.520 ;
        RECT 201.270 -29.780 201.530 -29.520 ;
        RECT 205.100 -29.780 205.360 -29.520 ;
        RECT 214.770 -29.780 215.030 -29.520 ;
        RECT 12.270 -30.560 12.530 -30.300 ;
        RECT 16.100 -30.560 16.360 -30.300 ;
        RECT 25.770 -30.560 26.030 -30.300 ;
        RECT 29.600 -30.560 29.860 -30.300 ;
        RECT 39.270 -30.560 39.530 -30.300 ;
        RECT 43.100 -30.560 43.360 -30.300 ;
        RECT 52.770 -30.560 53.030 -30.300 ;
        RECT 56.600 -30.560 56.860 -30.300 ;
        RECT 12.270 -33.390 12.530 -33.130 ;
        RECT 16.100 -33.390 16.360 -33.130 ;
        RECT 66.270 -30.560 66.530 -30.300 ;
        RECT 70.100 -30.560 70.360 -30.300 ;
        RECT 25.770 -33.390 26.030 -33.130 ;
        RECT 29.600 -33.390 29.860 -33.130 ;
        RECT 79.770 -30.560 80.030 -30.300 ;
        RECT 83.600 -30.560 83.860 -30.300 ;
        RECT 39.270 -33.390 39.530 -33.130 ;
        RECT 43.100 -33.390 43.360 -33.130 ;
        RECT 93.270 -30.560 93.530 -30.300 ;
        RECT 97.100 -30.560 97.360 -30.300 ;
        RECT 52.770 -33.390 53.030 -33.130 ;
        RECT 56.600 -33.390 56.860 -33.130 ;
        RECT 106.770 -30.560 107.030 -30.300 ;
        RECT 110.600 -30.560 110.860 -30.300 ;
        RECT 66.270 -33.390 66.530 -33.130 ;
        RECT 70.100 -33.390 70.360 -33.130 ;
        RECT 120.270 -30.560 120.530 -30.300 ;
        RECT 124.100 -30.560 124.360 -30.300 ;
        RECT 79.770 -33.390 80.030 -33.130 ;
        RECT 83.600 -33.390 83.860 -33.130 ;
        RECT 133.770 -30.560 134.030 -30.300 ;
        RECT 137.600 -30.560 137.860 -30.300 ;
        RECT 93.270 -33.390 93.530 -33.130 ;
        RECT 97.100 -33.390 97.360 -33.130 ;
        RECT 147.270 -30.560 147.530 -30.300 ;
        RECT 151.100 -30.560 151.360 -30.300 ;
        RECT 106.770 -33.390 107.030 -33.130 ;
        RECT 110.600 -33.390 110.860 -33.130 ;
        RECT 160.770 -30.560 161.030 -30.300 ;
        RECT 164.600 -30.560 164.860 -30.300 ;
        RECT 120.270 -33.390 120.530 -33.130 ;
        RECT 124.100 -33.390 124.360 -33.130 ;
        RECT 174.270 -30.560 174.530 -30.300 ;
        RECT 178.100 -30.560 178.360 -30.300 ;
        RECT 133.770 -33.390 134.030 -33.130 ;
        RECT 137.600 -33.390 137.860 -33.130 ;
        RECT 187.770 -30.560 188.030 -30.300 ;
        RECT 191.600 -30.560 191.860 -30.300 ;
        RECT 147.270 -33.390 147.530 -33.130 ;
        RECT 151.100 -33.390 151.360 -33.130 ;
        RECT 201.270 -30.560 201.530 -30.300 ;
        RECT 205.100 -30.560 205.360 -30.300 ;
        RECT 160.770 -33.390 161.030 -33.130 ;
        RECT 164.600 -33.390 164.860 -33.130 ;
        RECT 214.770 -30.560 215.030 -30.300 ;
        RECT 174.270 -33.390 174.530 -33.130 ;
        RECT 178.100 -33.390 178.360 -33.130 ;
        RECT 187.770 -33.390 188.030 -33.130 ;
        RECT 191.600 -33.390 191.860 -33.130 ;
        RECT 201.270 -33.390 201.530 -33.130 ;
        RECT 205.100 -33.390 205.360 -33.130 ;
        RECT 214.770 -33.390 215.030 -33.130 ;
        RECT 12.270 -34.170 12.530 -33.910 ;
        RECT 16.100 -34.170 16.360 -33.910 ;
        RECT 25.770 -34.170 26.030 -33.910 ;
        RECT 29.600 -34.170 29.860 -33.910 ;
        RECT 39.270 -34.170 39.530 -33.910 ;
        RECT 43.100 -34.170 43.360 -33.910 ;
        RECT 52.770 -34.170 53.030 -33.910 ;
        RECT 56.600 -34.170 56.860 -33.910 ;
        RECT 12.270 -37.000 12.530 -36.740 ;
        RECT 16.100 -37.000 16.360 -36.740 ;
        RECT 66.270 -34.170 66.530 -33.910 ;
        RECT 70.100 -34.170 70.360 -33.910 ;
        RECT 25.770 -37.000 26.030 -36.740 ;
        RECT 29.600 -37.000 29.860 -36.740 ;
        RECT 79.770 -34.170 80.030 -33.910 ;
        RECT 83.600 -34.170 83.860 -33.910 ;
        RECT 39.270 -37.000 39.530 -36.740 ;
        RECT 43.100 -37.000 43.360 -36.740 ;
        RECT 93.270 -34.170 93.530 -33.910 ;
        RECT 97.100 -34.170 97.360 -33.910 ;
        RECT 52.770 -37.000 53.030 -36.740 ;
        RECT 56.600 -37.000 56.860 -36.740 ;
        RECT 106.770 -34.170 107.030 -33.910 ;
        RECT 110.600 -34.170 110.860 -33.910 ;
        RECT 66.270 -37.000 66.530 -36.740 ;
        RECT 70.100 -37.000 70.360 -36.740 ;
        RECT 120.270 -34.170 120.530 -33.910 ;
        RECT 124.100 -34.170 124.360 -33.910 ;
        RECT 79.770 -37.000 80.030 -36.740 ;
        RECT 83.600 -37.000 83.860 -36.740 ;
        RECT 133.770 -34.170 134.030 -33.910 ;
        RECT 137.600 -34.170 137.860 -33.910 ;
        RECT 93.270 -37.000 93.530 -36.740 ;
        RECT 97.100 -37.000 97.360 -36.740 ;
        RECT 147.270 -34.170 147.530 -33.910 ;
        RECT 151.100 -34.170 151.360 -33.910 ;
        RECT 106.770 -37.000 107.030 -36.740 ;
        RECT 110.600 -37.000 110.860 -36.740 ;
        RECT 160.770 -34.170 161.030 -33.910 ;
        RECT 164.600 -34.170 164.860 -33.910 ;
        RECT 120.270 -37.000 120.530 -36.740 ;
        RECT 124.100 -37.000 124.360 -36.740 ;
        RECT 174.270 -34.170 174.530 -33.910 ;
        RECT 178.100 -34.170 178.360 -33.910 ;
        RECT 133.770 -37.000 134.030 -36.740 ;
        RECT 137.600 -37.000 137.860 -36.740 ;
        RECT 187.770 -34.170 188.030 -33.910 ;
        RECT 191.600 -34.170 191.860 -33.910 ;
        RECT 147.270 -37.000 147.530 -36.740 ;
        RECT 151.100 -37.000 151.360 -36.740 ;
        RECT 201.270 -34.170 201.530 -33.910 ;
        RECT 205.100 -34.170 205.360 -33.910 ;
        RECT 160.770 -37.000 161.030 -36.740 ;
        RECT 164.600 -37.000 164.860 -36.740 ;
        RECT 214.770 -34.170 215.030 -33.910 ;
        RECT 174.270 -37.000 174.530 -36.740 ;
        RECT 178.100 -37.000 178.360 -36.740 ;
        RECT 187.770 -37.000 188.030 -36.740 ;
        RECT 191.600 -37.000 191.860 -36.740 ;
        RECT 201.270 -37.000 201.530 -36.740 ;
        RECT 205.100 -37.000 205.360 -36.740 ;
        RECT 214.770 -37.000 215.030 -36.740 ;
        RECT 12.270 -37.780 12.530 -37.520 ;
        RECT 16.100 -37.780 16.360 -37.520 ;
        RECT 25.770 -37.780 26.030 -37.520 ;
        RECT 29.600 -37.780 29.860 -37.520 ;
        RECT 39.270 -37.780 39.530 -37.520 ;
        RECT 43.100 -37.780 43.360 -37.520 ;
        RECT 52.770 -37.780 53.030 -37.520 ;
        RECT 56.600 -37.780 56.860 -37.520 ;
        RECT 12.270 -40.610 12.530 -40.350 ;
        RECT 16.100 -40.610 16.360 -40.350 ;
        RECT 66.270 -37.780 66.530 -37.520 ;
        RECT 70.100 -37.780 70.360 -37.520 ;
        RECT 25.770 -40.610 26.030 -40.350 ;
        RECT 29.600 -40.610 29.860 -40.350 ;
        RECT 79.770 -37.780 80.030 -37.520 ;
        RECT 83.600 -37.780 83.860 -37.520 ;
        RECT 39.270 -40.610 39.530 -40.350 ;
        RECT 43.100 -40.610 43.360 -40.350 ;
        RECT 93.270 -37.780 93.530 -37.520 ;
        RECT 97.100 -37.780 97.360 -37.520 ;
        RECT 52.770 -40.610 53.030 -40.350 ;
        RECT 56.600 -40.610 56.860 -40.350 ;
        RECT 106.770 -37.780 107.030 -37.520 ;
        RECT 110.600 -37.780 110.860 -37.520 ;
        RECT 66.270 -40.610 66.530 -40.350 ;
        RECT 70.100 -40.610 70.360 -40.350 ;
        RECT 120.270 -37.780 120.530 -37.520 ;
        RECT 124.100 -37.780 124.360 -37.520 ;
        RECT 79.770 -40.610 80.030 -40.350 ;
        RECT 83.600 -40.610 83.860 -40.350 ;
        RECT 133.770 -37.780 134.030 -37.520 ;
        RECT 137.600 -37.780 137.860 -37.520 ;
        RECT 93.270 -40.610 93.530 -40.350 ;
        RECT 97.100 -40.610 97.360 -40.350 ;
        RECT 147.270 -37.780 147.530 -37.520 ;
        RECT 151.100 -37.780 151.360 -37.520 ;
        RECT 106.770 -40.610 107.030 -40.350 ;
        RECT 110.600 -40.610 110.860 -40.350 ;
        RECT 160.770 -37.780 161.030 -37.520 ;
        RECT 164.600 -37.780 164.860 -37.520 ;
        RECT 120.270 -40.610 120.530 -40.350 ;
        RECT 124.100 -40.610 124.360 -40.350 ;
        RECT 174.270 -37.780 174.530 -37.520 ;
        RECT 178.100 -37.780 178.360 -37.520 ;
        RECT 133.770 -40.610 134.030 -40.350 ;
        RECT 137.600 -40.610 137.860 -40.350 ;
        RECT 187.770 -37.780 188.030 -37.520 ;
        RECT 191.600 -37.780 191.860 -37.520 ;
        RECT 147.270 -40.610 147.530 -40.350 ;
        RECT 151.100 -40.610 151.360 -40.350 ;
        RECT 201.270 -37.780 201.530 -37.520 ;
        RECT 205.100 -37.780 205.360 -37.520 ;
        RECT 160.770 -40.610 161.030 -40.350 ;
        RECT 164.600 -40.610 164.860 -40.350 ;
        RECT 214.770 -37.780 215.030 -37.520 ;
        RECT 174.270 -40.610 174.530 -40.350 ;
        RECT 178.100 -40.610 178.360 -40.350 ;
        RECT 187.770 -40.610 188.030 -40.350 ;
        RECT 191.600 -40.610 191.860 -40.350 ;
        RECT 201.270 -40.610 201.530 -40.350 ;
        RECT 205.100 -40.610 205.360 -40.350 ;
        RECT 214.770 -40.610 215.030 -40.350 ;
      LAYER met1 ;
        RECT 9.180 -41.220 9.770 17.240 ;
        RECT 12.060 -41.200 12.630 17.220 ;
        RECT 16.000 -41.200 16.570 17.220 ;
        RECT 18.860 -41.220 19.450 17.240 ;
        RECT 22.680 -41.220 23.270 17.240 ;
        RECT 25.560 -41.200 26.130 17.220 ;
        RECT 29.500 -41.200 30.070 17.220 ;
        RECT 32.360 -41.220 32.950 17.240 ;
        RECT 36.180 -41.220 36.770 17.240 ;
        RECT 39.060 -41.200 39.630 17.220 ;
        RECT 43.000 -41.200 43.570 17.220 ;
        RECT 45.860 -41.220 46.450 17.240 ;
        RECT 49.680 -41.220 50.270 17.240 ;
        RECT 52.560 -41.200 53.130 17.220 ;
        RECT 56.500 -41.200 57.070 17.220 ;
        RECT 59.360 -41.220 59.950 17.240 ;
        RECT 63.180 -41.220 63.770 17.240 ;
        RECT 66.060 -41.200 66.630 17.220 ;
        RECT 70.000 -41.200 70.570 17.220 ;
        RECT 72.860 -41.220 73.450 17.240 ;
        RECT 76.680 -41.220 77.270 17.240 ;
        RECT 79.560 -41.200 80.130 17.220 ;
        RECT 83.500 -41.200 84.070 17.220 ;
        RECT 86.360 -41.220 86.950 17.240 ;
        RECT 90.180 -41.220 90.770 17.240 ;
        RECT 93.060 -41.200 93.630 17.220 ;
        RECT 97.000 -41.200 97.570 17.220 ;
        RECT 99.860 -41.220 100.450 17.240 ;
        RECT 103.680 -41.220 104.270 17.240 ;
        RECT 106.560 -41.200 107.130 17.220 ;
        RECT 110.500 -41.200 111.070 17.220 ;
        RECT 113.360 -41.220 113.950 17.240 ;
        RECT 117.180 -41.220 117.770 17.240 ;
        RECT 120.060 -41.200 120.630 17.220 ;
        RECT 124.000 -41.200 124.570 17.220 ;
        RECT 126.860 -41.220 127.450 17.240 ;
        RECT 130.680 -41.220 131.270 17.240 ;
        RECT 133.560 -41.200 134.130 17.220 ;
        RECT 137.500 -41.200 138.070 17.220 ;
        RECT 140.360 -41.220 140.950 17.240 ;
        RECT 144.180 -41.220 144.770 17.240 ;
        RECT 147.060 -41.200 147.630 17.220 ;
        RECT 151.000 -41.200 151.570 17.220 ;
        RECT 153.860 -41.220 154.450 17.240 ;
        RECT 157.680 -41.220 158.270 17.240 ;
        RECT 160.560 -41.200 161.130 17.220 ;
        RECT 164.500 -41.200 165.070 17.220 ;
        RECT 167.360 -41.220 167.950 17.240 ;
        RECT 171.180 -41.220 171.770 17.240 ;
        RECT 174.060 -41.200 174.630 17.220 ;
        RECT 178.000 -41.200 178.570 17.220 ;
        RECT 180.860 -41.220 181.450 17.240 ;
        RECT 184.680 -41.220 185.270 17.240 ;
        RECT 187.560 -41.200 188.130 17.220 ;
        RECT 191.500 -41.200 192.070 17.220 ;
        RECT 194.360 -41.220 194.950 17.240 ;
        RECT 198.180 -41.220 198.770 17.240 ;
        RECT 201.060 -41.200 201.630 17.220 ;
        RECT 205.000 -41.200 205.570 17.220 ;
        RECT 207.860 -41.220 208.450 17.240 ;
        RECT 211.680 -41.220 212.270 17.240 ;
        RECT 214.560 -41.200 215.130 17.220 ;
      LAYER via ;
        RECT 9.360 15.140 9.620 15.400 ;
        RECT 9.360 14.770 9.620 15.030 ;
        RECT 9.360 11.530 9.620 11.790 ;
        RECT 9.360 11.160 9.620 11.420 ;
        RECT 9.360 7.920 9.620 8.180 ;
        RECT 9.360 7.550 9.620 7.810 ;
        RECT 9.360 4.310 9.620 4.570 ;
        RECT 9.360 3.940 9.620 4.200 ;
        RECT 9.360 0.700 9.620 0.960 ;
        RECT 9.360 0.330 9.620 0.590 ;
        RECT 9.360 -2.910 9.620 -2.650 ;
        RECT 9.360 -3.280 9.620 -3.020 ;
        RECT 9.360 -6.520 9.620 -6.260 ;
        RECT 9.360 -6.890 9.620 -6.630 ;
        RECT 9.360 -10.130 9.620 -9.870 ;
        RECT 9.360 -10.500 9.620 -10.240 ;
        RECT 9.360 -13.740 9.620 -13.480 ;
        RECT 9.360 -14.110 9.620 -13.850 ;
        RECT 9.360 -17.350 9.620 -17.090 ;
        RECT 9.360 -17.720 9.620 -17.460 ;
        RECT 9.360 -20.960 9.620 -20.700 ;
        RECT 9.360 -21.330 9.620 -21.070 ;
        RECT 9.360 -24.570 9.620 -24.310 ;
        RECT 9.360 -24.940 9.620 -24.680 ;
        RECT 9.360 -28.180 9.620 -27.920 ;
        RECT 9.360 -28.550 9.620 -28.290 ;
        RECT 9.360 -31.790 9.620 -31.530 ;
        RECT 9.360 -32.160 9.620 -31.900 ;
        RECT 9.360 -35.400 9.620 -35.140 ;
        RECT 9.360 -35.770 9.620 -35.510 ;
        RECT 9.360 -39.010 9.620 -38.750 ;
        RECT 9.360 -39.380 9.620 -39.120 ;
        RECT 12.220 15.130 12.480 15.390 ;
        RECT 12.220 14.780 12.480 15.040 ;
        RECT 12.220 11.520 12.480 11.780 ;
        RECT 12.220 11.170 12.480 11.430 ;
        RECT 12.220 7.910 12.480 8.170 ;
        RECT 12.220 7.560 12.480 7.820 ;
        RECT 12.220 4.300 12.480 4.560 ;
        RECT 12.220 3.950 12.480 4.210 ;
        RECT 12.220 0.690 12.480 0.950 ;
        RECT 12.220 0.340 12.480 0.600 ;
        RECT 12.220 -2.920 12.480 -2.660 ;
        RECT 12.220 -3.270 12.480 -3.010 ;
        RECT 12.220 -6.530 12.480 -6.270 ;
        RECT 12.220 -6.880 12.480 -6.620 ;
        RECT 12.220 -10.140 12.480 -9.880 ;
        RECT 12.220 -10.490 12.480 -10.230 ;
        RECT 12.220 -13.750 12.480 -13.490 ;
        RECT 12.220 -14.100 12.480 -13.840 ;
        RECT 12.220 -17.360 12.480 -17.100 ;
        RECT 12.220 -17.710 12.480 -17.450 ;
        RECT 12.220 -20.970 12.480 -20.710 ;
        RECT 12.220 -21.320 12.480 -21.060 ;
        RECT 12.220 -24.580 12.480 -24.320 ;
        RECT 12.220 -24.930 12.480 -24.670 ;
        RECT 12.220 -28.190 12.480 -27.930 ;
        RECT 12.220 -28.540 12.480 -28.280 ;
        RECT 12.220 -31.800 12.480 -31.540 ;
        RECT 12.220 -32.150 12.480 -31.890 ;
        RECT 12.220 -35.410 12.480 -35.150 ;
        RECT 12.220 -35.760 12.480 -35.500 ;
        RECT 12.220 -39.020 12.480 -38.760 ;
        RECT 12.220 -39.370 12.480 -39.110 ;
        RECT 16.150 15.130 16.410 15.390 ;
        RECT 16.150 14.780 16.410 15.040 ;
        RECT 16.150 11.520 16.410 11.780 ;
        RECT 16.150 11.170 16.410 11.430 ;
        RECT 16.150 7.910 16.410 8.170 ;
        RECT 16.150 7.560 16.410 7.820 ;
        RECT 16.150 4.300 16.410 4.560 ;
        RECT 16.150 3.950 16.410 4.210 ;
        RECT 16.150 0.690 16.410 0.950 ;
        RECT 16.150 0.340 16.410 0.600 ;
        RECT 16.150 -2.920 16.410 -2.660 ;
        RECT 16.150 -3.270 16.410 -3.010 ;
        RECT 16.150 -6.530 16.410 -6.270 ;
        RECT 16.150 -6.880 16.410 -6.620 ;
        RECT 16.150 -10.140 16.410 -9.880 ;
        RECT 16.150 -10.490 16.410 -10.230 ;
        RECT 16.150 -13.750 16.410 -13.490 ;
        RECT 16.150 -14.100 16.410 -13.840 ;
        RECT 16.150 -17.360 16.410 -17.100 ;
        RECT 16.150 -17.710 16.410 -17.450 ;
        RECT 16.150 -20.970 16.410 -20.710 ;
        RECT 16.150 -21.320 16.410 -21.060 ;
        RECT 16.150 -24.580 16.410 -24.320 ;
        RECT 16.150 -24.930 16.410 -24.670 ;
        RECT 16.150 -28.190 16.410 -27.930 ;
        RECT 16.150 -28.540 16.410 -28.280 ;
        RECT 16.150 -31.800 16.410 -31.540 ;
        RECT 16.150 -32.150 16.410 -31.890 ;
        RECT 16.150 -35.410 16.410 -35.150 ;
        RECT 16.150 -35.760 16.410 -35.500 ;
        RECT 16.150 -39.020 16.410 -38.760 ;
        RECT 16.150 -39.370 16.410 -39.110 ;
        RECT 19.010 15.140 19.270 15.400 ;
        RECT 19.010 14.770 19.270 15.030 ;
        RECT 19.010 11.530 19.270 11.790 ;
        RECT 19.010 11.160 19.270 11.420 ;
        RECT 19.010 7.920 19.270 8.180 ;
        RECT 19.010 7.550 19.270 7.810 ;
        RECT 19.010 4.310 19.270 4.570 ;
        RECT 19.010 3.940 19.270 4.200 ;
        RECT 19.010 0.700 19.270 0.960 ;
        RECT 19.010 0.330 19.270 0.590 ;
        RECT 19.010 -2.910 19.270 -2.650 ;
        RECT 19.010 -3.280 19.270 -3.020 ;
        RECT 19.010 -6.520 19.270 -6.260 ;
        RECT 19.010 -6.890 19.270 -6.630 ;
        RECT 19.010 -10.130 19.270 -9.870 ;
        RECT 19.010 -10.500 19.270 -10.240 ;
        RECT 19.010 -13.740 19.270 -13.480 ;
        RECT 19.010 -14.110 19.270 -13.850 ;
        RECT 19.010 -17.350 19.270 -17.090 ;
        RECT 19.010 -17.720 19.270 -17.460 ;
        RECT 19.010 -20.960 19.270 -20.700 ;
        RECT 19.010 -21.330 19.270 -21.070 ;
        RECT 19.010 -24.570 19.270 -24.310 ;
        RECT 19.010 -24.940 19.270 -24.680 ;
        RECT 19.010 -28.180 19.270 -27.920 ;
        RECT 19.010 -28.550 19.270 -28.290 ;
        RECT 19.010 -31.790 19.270 -31.530 ;
        RECT 19.010 -32.160 19.270 -31.900 ;
        RECT 19.010 -35.400 19.270 -35.140 ;
        RECT 19.010 -35.770 19.270 -35.510 ;
        RECT 19.010 -39.010 19.270 -38.750 ;
        RECT 19.010 -39.380 19.270 -39.120 ;
        RECT 22.860 15.140 23.120 15.400 ;
        RECT 22.860 14.770 23.120 15.030 ;
        RECT 22.860 11.530 23.120 11.790 ;
        RECT 22.860 11.160 23.120 11.420 ;
        RECT 22.860 7.920 23.120 8.180 ;
        RECT 22.860 7.550 23.120 7.810 ;
        RECT 22.860 4.310 23.120 4.570 ;
        RECT 22.860 3.940 23.120 4.200 ;
        RECT 22.860 0.700 23.120 0.960 ;
        RECT 22.860 0.330 23.120 0.590 ;
        RECT 22.860 -2.910 23.120 -2.650 ;
        RECT 22.860 -3.280 23.120 -3.020 ;
        RECT 22.860 -6.520 23.120 -6.260 ;
        RECT 22.860 -6.890 23.120 -6.630 ;
        RECT 22.860 -10.130 23.120 -9.870 ;
        RECT 22.860 -10.500 23.120 -10.240 ;
        RECT 22.860 -13.740 23.120 -13.480 ;
        RECT 22.860 -14.110 23.120 -13.850 ;
        RECT 22.860 -17.350 23.120 -17.090 ;
        RECT 22.860 -17.720 23.120 -17.460 ;
        RECT 22.860 -20.960 23.120 -20.700 ;
        RECT 22.860 -21.330 23.120 -21.070 ;
        RECT 22.860 -24.570 23.120 -24.310 ;
        RECT 22.860 -24.940 23.120 -24.680 ;
        RECT 22.860 -28.180 23.120 -27.920 ;
        RECT 22.860 -28.550 23.120 -28.290 ;
        RECT 22.860 -31.790 23.120 -31.530 ;
        RECT 22.860 -32.160 23.120 -31.900 ;
        RECT 22.860 -35.400 23.120 -35.140 ;
        RECT 22.860 -35.770 23.120 -35.510 ;
        RECT 22.860 -39.010 23.120 -38.750 ;
        RECT 22.860 -39.380 23.120 -39.120 ;
        RECT 25.720 15.130 25.980 15.390 ;
        RECT 25.720 14.780 25.980 15.040 ;
        RECT 25.720 11.520 25.980 11.780 ;
        RECT 25.720 11.170 25.980 11.430 ;
        RECT 25.720 7.910 25.980 8.170 ;
        RECT 25.720 7.560 25.980 7.820 ;
        RECT 25.720 4.300 25.980 4.560 ;
        RECT 25.720 3.950 25.980 4.210 ;
        RECT 25.720 0.690 25.980 0.950 ;
        RECT 25.720 0.340 25.980 0.600 ;
        RECT 25.720 -2.920 25.980 -2.660 ;
        RECT 25.720 -3.270 25.980 -3.010 ;
        RECT 25.720 -6.530 25.980 -6.270 ;
        RECT 25.720 -6.880 25.980 -6.620 ;
        RECT 25.720 -10.140 25.980 -9.880 ;
        RECT 25.720 -10.490 25.980 -10.230 ;
        RECT 25.720 -13.750 25.980 -13.490 ;
        RECT 25.720 -14.100 25.980 -13.840 ;
        RECT 25.720 -17.360 25.980 -17.100 ;
        RECT 25.720 -17.710 25.980 -17.450 ;
        RECT 25.720 -20.970 25.980 -20.710 ;
        RECT 25.720 -21.320 25.980 -21.060 ;
        RECT 25.720 -24.580 25.980 -24.320 ;
        RECT 25.720 -24.930 25.980 -24.670 ;
        RECT 25.720 -28.190 25.980 -27.930 ;
        RECT 25.720 -28.540 25.980 -28.280 ;
        RECT 25.720 -31.800 25.980 -31.540 ;
        RECT 25.720 -32.150 25.980 -31.890 ;
        RECT 25.720 -35.410 25.980 -35.150 ;
        RECT 25.720 -35.760 25.980 -35.500 ;
        RECT 25.720 -39.020 25.980 -38.760 ;
        RECT 25.720 -39.370 25.980 -39.110 ;
        RECT 29.650 15.130 29.910 15.390 ;
        RECT 29.650 14.780 29.910 15.040 ;
        RECT 29.650 11.520 29.910 11.780 ;
        RECT 29.650 11.170 29.910 11.430 ;
        RECT 29.650 7.910 29.910 8.170 ;
        RECT 29.650 7.560 29.910 7.820 ;
        RECT 29.650 4.300 29.910 4.560 ;
        RECT 29.650 3.950 29.910 4.210 ;
        RECT 29.650 0.690 29.910 0.950 ;
        RECT 29.650 0.340 29.910 0.600 ;
        RECT 29.650 -2.920 29.910 -2.660 ;
        RECT 29.650 -3.270 29.910 -3.010 ;
        RECT 29.650 -6.530 29.910 -6.270 ;
        RECT 29.650 -6.880 29.910 -6.620 ;
        RECT 29.650 -10.140 29.910 -9.880 ;
        RECT 29.650 -10.490 29.910 -10.230 ;
        RECT 29.650 -13.750 29.910 -13.490 ;
        RECT 29.650 -14.100 29.910 -13.840 ;
        RECT 29.650 -17.360 29.910 -17.100 ;
        RECT 29.650 -17.710 29.910 -17.450 ;
        RECT 29.650 -20.970 29.910 -20.710 ;
        RECT 29.650 -21.320 29.910 -21.060 ;
        RECT 29.650 -24.580 29.910 -24.320 ;
        RECT 29.650 -24.930 29.910 -24.670 ;
        RECT 29.650 -28.190 29.910 -27.930 ;
        RECT 29.650 -28.540 29.910 -28.280 ;
        RECT 29.650 -31.800 29.910 -31.540 ;
        RECT 29.650 -32.150 29.910 -31.890 ;
        RECT 29.650 -35.410 29.910 -35.150 ;
        RECT 29.650 -35.760 29.910 -35.500 ;
        RECT 29.650 -39.020 29.910 -38.760 ;
        RECT 29.650 -39.370 29.910 -39.110 ;
        RECT 32.510 15.140 32.770 15.400 ;
        RECT 32.510 14.770 32.770 15.030 ;
        RECT 32.510 11.530 32.770 11.790 ;
        RECT 32.510 11.160 32.770 11.420 ;
        RECT 32.510 7.920 32.770 8.180 ;
        RECT 32.510 7.550 32.770 7.810 ;
        RECT 32.510 4.310 32.770 4.570 ;
        RECT 32.510 3.940 32.770 4.200 ;
        RECT 32.510 0.700 32.770 0.960 ;
        RECT 32.510 0.330 32.770 0.590 ;
        RECT 32.510 -2.910 32.770 -2.650 ;
        RECT 32.510 -3.280 32.770 -3.020 ;
        RECT 32.510 -6.520 32.770 -6.260 ;
        RECT 32.510 -6.890 32.770 -6.630 ;
        RECT 32.510 -10.130 32.770 -9.870 ;
        RECT 32.510 -10.500 32.770 -10.240 ;
        RECT 32.510 -13.740 32.770 -13.480 ;
        RECT 32.510 -14.110 32.770 -13.850 ;
        RECT 32.510 -17.350 32.770 -17.090 ;
        RECT 32.510 -17.720 32.770 -17.460 ;
        RECT 32.510 -20.960 32.770 -20.700 ;
        RECT 32.510 -21.330 32.770 -21.070 ;
        RECT 32.510 -24.570 32.770 -24.310 ;
        RECT 32.510 -24.940 32.770 -24.680 ;
        RECT 32.510 -28.180 32.770 -27.920 ;
        RECT 32.510 -28.550 32.770 -28.290 ;
        RECT 32.510 -31.790 32.770 -31.530 ;
        RECT 32.510 -32.160 32.770 -31.900 ;
        RECT 32.510 -35.400 32.770 -35.140 ;
        RECT 32.510 -35.770 32.770 -35.510 ;
        RECT 32.510 -39.010 32.770 -38.750 ;
        RECT 32.510 -39.380 32.770 -39.120 ;
        RECT 36.360 15.140 36.620 15.400 ;
        RECT 36.360 14.770 36.620 15.030 ;
        RECT 36.360 11.530 36.620 11.790 ;
        RECT 36.360 11.160 36.620 11.420 ;
        RECT 36.360 7.920 36.620 8.180 ;
        RECT 36.360 7.550 36.620 7.810 ;
        RECT 36.360 4.310 36.620 4.570 ;
        RECT 36.360 3.940 36.620 4.200 ;
        RECT 36.360 0.700 36.620 0.960 ;
        RECT 36.360 0.330 36.620 0.590 ;
        RECT 36.360 -2.910 36.620 -2.650 ;
        RECT 36.360 -3.280 36.620 -3.020 ;
        RECT 36.360 -6.520 36.620 -6.260 ;
        RECT 36.360 -6.890 36.620 -6.630 ;
        RECT 36.360 -10.130 36.620 -9.870 ;
        RECT 36.360 -10.500 36.620 -10.240 ;
        RECT 36.360 -13.740 36.620 -13.480 ;
        RECT 36.360 -14.110 36.620 -13.850 ;
        RECT 36.360 -17.350 36.620 -17.090 ;
        RECT 36.360 -17.720 36.620 -17.460 ;
        RECT 36.360 -20.960 36.620 -20.700 ;
        RECT 36.360 -21.330 36.620 -21.070 ;
        RECT 36.360 -24.570 36.620 -24.310 ;
        RECT 36.360 -24.940 36.620 -24.680 ;
        RECT 36.360 -28.180 36.620 -27.920 ;
        RECT 36.360 -28.550 36.620 -28.290 ;
        RECT 36.360 -31.790 36.620 -31.530 ;
        RECT 36.360 -32.160 36.620 -31.900 ;
        RECT 36.360 -35.400 36.620 -35.140 ;
        RECT 36.360 -35.770 36.620 -35.510 ;
        RECT 36.360 -39.010 36.620 -38.750 ;
        RECT 36.360 -39.380 36.620 -39.120 ;
        RECT 39.220 15.130 39.480 15.390 ;
        RECT 39.220 14.780 39.480 15.040 ;
        RECT 39.220 11.520 39.480 11.780 ;
        RECT 39.220 11.170 39.480 11.430 ;
        RECT 39.220 7.910 39.480 8.170 ;
        RECT 39.220 7.560 39.480 7.820 ;
        RECT 39.220 4.300 39.480 4.560 ;
        RECT 39.220 3.950 39.480 4.210 ;
        RECT 39.220 0.690 39.480 0.950 ;
        RECT 39.220 0.340 39.480 0.600 ;
        RECT 39.220 -2.920 39.480 -2.660 ;
        RECT 39.220 -3.270 39.480 -3.010 ;
        RECT 39.220 -6.530 39.480 -6.270 ;
        RECT 39.220 -6.880 39.480 -6.620 ;
        RECT 39.220 -10.140 39.480 -9.880 ;
        RECT 39.220 -10.490 39.480 -10.230 ;
        RECT 39.220 -13.750 39.480 -13.490 ;
        RECT 39.220 -14.100 39.480 -13.840 ;
        RECT 39.220 -17.360 39.480 -17.100 ;
        RECT 39.220 -17.710 39.480 -17.450 ;
        RECT 39.220 -20.970 39.480 -20.710 ;
        RECT 39.220 -21.320 39.480 -21.060 ;
        RECT 39.220 -24.580 39.480 -24.320 ;
        RECT 39.220 -24.930 39.480 -24.670 ;
        RECT 39.220 -28.190 39.480 -27.930 ;
        RECT 39.220 -28.540 39.480 -28.280 ;
        RECT 39.220 -31.800 39.480 -31.540 ;
        RECT 39.220 -32.150 39.480 -31.890 ;
        RECT 39.220 -35.410 39.480 -35.150 ;
        RECT 39.220 -35.760 39.480 -35.500 ;
        RECT 39.220 -39.020 39.480 -38.760 ;
        RECT 39.220 -39.370 39.480 -39.110 ;
        RECT 43.150 15.130 43.410 15.390 ;
        RECT 43.150 14.780 43.410 15.040 ;
        RECT 43.150 11.520 43.410 11.780 ;
        RECT 43.150 11.170 43.410 11.430 ;
        RECT 43.150 7.910 43.410 8.170 ;
        RECT 43.150 7.560 43.410 7.820 ;
        RECT 43.150 4.300 43.410 4.560 ;
        RECT 43.150 3.950 43.410 4.210 ;
        RECT 43.150 0.690 43.410 0.950 ;
        RECT 43.150 0.340 43.410 0.600 ;
        RECT 43.150 -2.920 43.410 -2.660 ;
        RECT 43.150 -3.270 43.410 -3.010 ;
        RECT 43.150 -6.530 43.410 -6.270 ;
        RECT 43.150 -6.880 43.410 -6.620 ;
        RECT 43.150 -10.140 43.410 -9.880 ;
        RECT 43.150 -10.490 43.410 -10.230 ;
        RECT 43.150 -13.750 43.410 -13.490 ;
        RECT 43.150 -14.100 43.410 -13.840 ;
        RECT 43.150 -17.360 43.410 -17.100 ;
        RECT 43.150 -17.710 43.410 -17.450 ;
        RECT 43.150 -20.970 43.410 -20.710 ;
        RECT 43.150 -21.320 43.410 -21.060 ;
        RECT 43.150 -24.580 43.410 -24.320 ;
        RECT 43.150 -24.930 43.410 -24.670 ;
        RECT 43.150 -28.190 43.410 -27.930 ;
        RECT 43.150 -28.540 43.410 -28.280 ;
        RECT 43.150 -31.800 43.410 -31.540 ;
        RECT 43.150 -32.150 43.410 -31.890 ;
        RECT 43.150 -35.410 43.410 -35.150 ;
        RECT 43.150 -35.760 43.410 -35.500 ;
        RECT 43.150 -39.020 43.410 -38.760 ;
        RECT 43.150 -39.370 43.410 -39.110 ;
        RECT 46.010 15.140 46.270 15.400 ;
        RECT 46.010 14.770 46.270 15.030 ;
        RECT 46.010 11.530 46.270 11.790 ;
        RECT 46.010 11.160 46.270 11.420 ;
        RECT 46.010 7.920 46.270 8.180 ;
        RECT 46.010 7.550 46.270 7.810 ;
        RECT 46.010 4.310 46.270 4.570 ;
        RECT 46.010 3.940 46.270 4.200 ;
        RECT 46.010 0.700 46.270 0.960 ;
        RECT 46.010 0.330 46.270 0.590 ;
        RECT 46.010 -2.910 46.270 -2.650 ;
        RECT 46.010 -3.280 46.270 -3.020 ;
        RECT 46.010 -6.520 46.270 -6.260 ;
        RECT 46.010 -6.890 46.270 -6.630 ;
        RECT 46.010 -10.130 46.270 -9.870 ;
        RECT 46.010 -10.500 46.270 -10.240 ;
        RECT 46.010 -13.740 46.270 -13.480 ;
        RECT 46.010 -14.110 46.270 -13.850 ;
        RECT 46.010 -17.350 46.270 -17.090 ;
        RECT 46.010 -17.720 46.270 -17.460 ;
        RECT 46.010 -20.960 46.270 -20.700 ;
        RECT 46.010 -21.330 46.270 -21.070 ;
        RECT 46.010 -24.570 46.270 -24.310 ;
        RECT 46.010 -24.940 46.270 -24.680 ;
        RECT 46.010 -28.180 46.270 -27.920 ;
        RECT 46.010 -28.550 46.270 -28.290 ;
        RECT 46.010 -31.790 46.270 -31.530 ;
        RECT 46.010 -32.160 46.270 -31.900 ;
        RECT 46.010 -35.400 46.270 -35.140 ;
        RECT 46.010 -35.770 46.270 -35.510 ;
        RECT 46.010 -39.010 46.270 -38.750 ;
        RECT 46.010 -39.380 46.270 -39.120 ;
        RECT 49.860 15.140 50.120 15.400 ;
        RECT 49.860 14.770 50.120 15.030 ;
        RECT 49.860 11.530 50.120 11.790 ;
        RECT 49.860 11.160 50.120 11.420 ;
        RECT 49.860 7.920 50.120 8.180 ;
        RECT 49.860 7.550 50.120 7.810 ;
        RECT 49.860 4.310 50.120 4.570 ;
        RECT 49.860 3.940 50.120 4.200 ;
        RECT 49.860 0.700 50.120 0.960 ;
        RECT 49.860 0.330 50.120 0.590 ;
        RECT 49.860 -2.910 50.120 -2.650 ;
        RECT 49.860 -3.280 50.120 -3.020 ;
        RECT 49.860 -6.520 50.120 -6.260 ;
        RECT 49.860 -6.890 50.120 -6.630 ;
        RECT 49.860 -10.130 50.120 -9.870 ;
        RECT 49.860 -10.500 50.120 -10.240 ;
        RECT 49.860 -13.740 50.120 -13.480 ;
        RECT 49.860 -14.110 50.120 -13.850 ;
        RECT 49.860 -17.350 50.120 -17.090 ;
        RECT 49.860 -17.720 50.120 -17.460 ;
        RECT 49.860 -20.960 50.120 -20.700 ;
        RECT 49.860 -21.330 50.120 -21.070 ;
        RECT 49.860 -24.570 50.120 -24.310 ;
        RECT 49.860 -24.940 50.120 -24.680 ;
        RECT 49.860 -28.180 50.120 -27.920 ;
        RECT 49.860 -28.550 50.120 -28.290 ;
        RECT 49.860 -31.790 50.120 -31.530 ;
        RECT 49.860 -32.160 50.120 -31.900 ;
        RECT 49.860 -35.400 50.120 -35.140 ;
        RECT 49.860 -35.770 50.120 -35.510 ;
        RECT 49.860 -39.010 50.120 -38.750 ;
        RECT 49.860 -39.380 50.120 -39.120 ;
        RECT 52.720 15.130 52.980 15.390 ;
        RECT 52.720 14.780 52.980 15.040 ;
        RECT 52.720 11.520 52.980 11.780 ;
        RECT 52.720 11.170 52.980 11.430 ;
        RECT 52.720 7.910 52.980 8.170 ;
        RECT 52.720 7.560 52.980 7.820 ;
        RECT 52.720 4.300 52.980 4.560 ;
        RECT 52.720 3.950 52.980 4.210 ;
        RECT 52.720 0.690 52.980 0.950 ;
        RECT 52.720 0.340 52.980 0.600 ;
        RECT 52.720 -2.920 52.980 -2.660 ;
        RECT 52.720 -3.270 52.980 -3.010 ;
        RECT 52.720 -6.530 52.980 -6.270 ;
        RECT 52.720 -6.880 52.980 -6.620 ;
        RECT 52.720 -10.140 52.980 -9.880 ;
        RECT 52.720 -10.490 52.980 -10.230 ;
        RECT 52.720 -13.750 52.980 -13.490 ;
        RECT 52.720 -14.100 52.980 -13.840 ;
        RECT 52.720 -17.360 52.980 -17.100 ;
        RECT 52.720 -17.710 52.980 -17.450 ;
        RECT 52.720 -20.970 52.980 -20.710 ;
        RECT 52.720 -21.320 52.980 -21.060 ;
        RECT 52.720 -24.580 52.980 -24.320 ;
        RECT 52.720 -24.930 52.980 -24.670 ;
        RECT 52.720 -28.190 52.980 -27.930 ;
        RECT 52.720 -28.540 52.980 -28.280 ;
        RECT 52.720 -31.800 52.980 -31.540 ;
        RECT 52.720 -32.150 52.980 -31.890 ;
        RECT 52.720 -35.410 52.980 -35.150 ;
        RECT 52.720 -35.760 52.980 -35.500 ;
        RECT 52.720 -39.020 52.980 -38.760 ;
        RECT 52.720 -39.370 52.980 -39.110 ;
        RECT 56.650 15.130 56.910 15.390 ;
        RECT 56.650 14.780 56.910 15.040 ;
        RECT 56.650 11.520 56.910 11.780 ;
        RECT 56.650 11.170 56.910 11.430 ;
        RECT 56.650 7.910 56.910 8.170 ;
        RECT 56.650 7.560 56.910 7.820 ;
        RECT 56.650 4.300 56.910 4.560 ;
        RECT 56.650 3.950 56.910 4.210 ;
        RECT 56.650 0.690 56.910 0.950 ;
        RECT 56.650 0.340 56.910 0.600 ;
        RECT 56.650 -2.920 56.910 -2.660 ;
        RECT 56.650 -3.270 56.910 -3.010 ;
        RECT 56.650 -6.530 56.910 -6.270 ;
        RECT 56.650 -6.880 56.910 -6.620 ;
        RECT 56.650 -10.140 56.910 -9.880 ;
        RECT 56.650 -10.490 56.910 -10.230 ;
        RECT 56.650 -13.750 56.910 -13.490 ;
        RECT 56.650 -14.100 56.910 -13.840 ;
        RECT 56.650 -17.360 56.910 -17.100 ;
        RECT 56.650 -17.710 56.910 -17.450 ;
        RECT 56.650 -20.970 56.910 -20.710 ;
        RECT 56.650 -21.320 56.910 -21.060 ;
        RECT 56.650 -24.580 56.910 -24.320 ;
        RECT 56.650 -24.930 56.910 -24.670 ;
        RECT 56.650 -28.190 56.910 -27.930 ;
        RECT 56.650 -28.540 56.910 -28.280 ;
        RECT 56.650 -31.800 56.910 -31.540 ;
        RECT 56.650 -32.150 56.910 -31.890 ;
        RECT 56.650 -35.410 56.910 -35.150 ;
        RECT 56.650 -35.760 56.910 -35.500 ;
        RECT 56.650 -39.020 56.910 -38.760 ;
        RECT 56.650 -39.370 56.910 -39.110 ;
        RECT 59.510 15.140 59.770 15.400 ;
        RECT 59.510 14.770 59.770 15.030 ;
        RECT 59.510 11.530 59.770 11.790 ;
        RECT 59.510 11.160 59.770 11.420 ;
        RECT 59.510 7.920 59.770 8.180 ;
        RECT 59.510 7.550 59.770 7.810 ;
        RECT 59.510 4.310 59.770 4.570 ;
        RECT 59.510 3.940 59.770 4.200 ;
        RECT 59.510 0.700 59.770 0.960 ;
        RECT 59.510 0.330 59.770 0.590 ;
        RECT 59.510 -2.910 59.770 -2.650 ;
        RECT 59.510 -3.280 59.770 -3.020 ;
        RECT 59.510 -6.520 59.770 -6.260 ;
        RECT 59.510 -6.890 59.770 -6.630 ;
        RECT 59.510 -10.130 59.770 -9.870 ;
        RECT 59.510 -10.500 59.770 -10.240 ;
        RECT 59.510 -13.740 59.770 -13.480 ;
        RECT 59.510 -14.110 59.770 -13.850 ;
        RECT 59.510 -17.350 59.770 -17.090 ;
        RECT 59.510 -17.720 59.770 -17.460 ;
        RECT 59.510 -20.960 59.770 -20.700 ;
        RECT 59.510 -21.330 59.770 -21.070 ;
        RECT 59.510 -24.570 59.770 -24.310 ;
        RECT 59.510 -24.940 59.770 -24.680 ;
        RECT 59.510 -28.180 59.770 -27.920 ;
        RECT 59.510 -28.550 59.770 -28.290 ;
        RECT 59.510 -31.790 59.770 -31.530 ;
        RECT 59.510 -32.160 59.770 -31.900 ;
        RECT 59.510 -35.400 59.770 -35.140 ;
        RECT 59.510 -35.770 59.770 -35.510 ;
        RECT 59.510 -39.010 59.770 -38.750 ;
        RECT 59.510 -39.380 59.770 -39.120 ;
        RECT 63.360 15.140 63.620 15.400 ;
        RECT 63.360 14.770 63.620 15.030 ;
        RECT 63.360 11.530 63.620 11.790 ;
        RECT 63.360 11.160 63.620 11.420 ;
        RECT 63.360 7.920 63.620 8.180 ;
        RECT 63.360 7.550 63.620 7.810 ;
        RECT 63.360 4.310 63.620 4.570 ;
        RECT 63.360 3.940 63.620 4.200 ;
        RECT 63.360 0.700 63.620 0.960 ;
        RECT 63.360 0.330 63.620 0.590 ;
        RECT 63.360 -2.910 63.620 -2.650 ;
        RECT 63.360 -3.280 63.620 -3.020 ;
        RECT 63.360 -6.520 63.620 -6.260 ;
        RECT 63.360 -6.890 63.620 -6.630 ;
        RECT 63.360 -10.130 63.620 -9.870 ;
        RECT 63.360 -10.500 63.620 -10.240 ;
        RECT 63.360 -13.740 63.620 -13.480 ;
        RECT 63.360 -14.110 63.620 -13.850 ;
        RECT 63.360 -17.350 63.620 -17.090 ;
        RECT 63.360 -17.720 63.620 -17.460 ;
        RECT 63.360 -20.960 63.620 -20.700 ;
        RECT 63.360 -21.330 63.620 -21.070 ;
        RECT 63.360 -24.570 63.620 -24.310 ;
        RECT 63.360 -24.940 63.620 -24.680 ;
        RECT 63.360 -28.180 63.620 -27.920 ;
        RECT 63.360 -28.550 63.620 -28.290 ;
        RECT 63.360 -31.790 63.620 -31.530 ;
        RECT 63.360 -32.160 63.620 -31.900 ;
        RECT 63.360 -35.400 63.620 -35.140 ;
        RECT 63.360 -35.770 63.620 -35.510 ;
        RECT 63.360 -39.010 63.620 -38.750 ;
        RECT 63.360 -39.380 63.620 -39.120 ;
        RECT 66.220 15.130 66.480 15.390 ;
        RECT 66.220 14.780 66.480 15.040 ;
        RECT 66.220 11.520 66.480 11.780 ;
        RECT 66.220 11.170 66.480 11.430 ;
        RECT 66.220 7.910 66.480 8.170 ;
        RECT 66.220 7.560 66.480 7.820 ;
        RECT 66.220 4.300 66.480 4.560 ;
        RECT 66.220 3.950 66.480 4.210 ;
        RECT 66.220 0.690 66.480 0.950 ;
        RECT 66.220 0.340 66.480 0.600 ;
        RECT 66.220 -2.920 66.480 -2.660 ;
        RECT 66.220 -3.270 66.480 -3.010 ;
        RECT 66.220 -6.530 66.480 -6.270 ;
        RECT 66.220 -6.880 66.480 -6.620 ;
        RECT 66.220 -10.140 66.480 -9.880 ;
        RECT 66.220 -10.490 66.480 -10.230 ;
        RECT 66.220 -13.750 66.480 -13.490 ;
        RECT 66.220 -14.100 66.480 -13.840 ;
        RECT 66.220 -17.360 66.480 -17.100 ;
        RECT 66.220 -17.710 66.480 -17.450 ;
        RECT 66.220 -20.970 66.480 -20.710 ;
        RECT 66.220 -21.320 66.480 -21.060 ;
        RECT 66.220 -24.580 66.480 -24.320 ;
        RECT 66.220 -24.930 66.480 -24.670 ;
        RECT 66.220 -28.190 66.480 -27.930 ;
        RECT 66.220 -28.540 66.480 -28.280 ;
        RECT 66.220 -31.800 66.480 -31.540 ;
        RECT 66.220 -32.150 66.480 -31.890 ;
        RECT 66.220 -35.410 66.480 -35.150 ;
        RECT 66.220 -35.760 66.480 -35.500 ;
        RECT 66.220 -39.020 66.480 -38.760 ;
        RECT 66.220 -39.370 66.480 -39.110 ;
        RECT 70.150 15.130 70.410 15.390 ;
        RECT 70.150 14.780 70.410 15.040 ;
        RECT 70.150 11.520 70.410 11.780 ;
        RECT 70.150 11.170 70.410 11.430 ;
        RECT 70.150 7.910 70.410 8.170 ;
        RECT 70.150 7.560 70.410 7.820 ;
        RECT 70.150 4.300 70.410 4.560 ;
        RECT 70.150 3.950 70.410 4.210 ;
        RECT 70.150 0.690 70.410 0.950 ;
        RECT 70.150 0.340 70.410 0.600 ;
        RECT 70.150 -2.920 70.410 -2.660 ;
        RECT 70.150 -3.270 70.410 -3.010 ;
        RECT 70.150 -6.530 70.410 -6.270 ;
        RECT 70.150 -6.880 70.410 -6.620 ;
        RECT 70.150 -10.140 70.410 -9.880 ;
        RECT 70.150 -10.490 70.410 -10.230 ;
        RECT 70.150 -13.750 70.410 -13.490 ;
        RECT 70.150 -14.100 70.410 -13.840 ;
        RECT 70.150 -17.360 70.410 -17.100 ;
        RECT 70.150 -17.710 70.410 -17.450 ;
        RECT 70.150 -20.970 70.410 -20.710 ;
        RECT 70.150 -21.320 70.410 -21.060 ;
        RECT 70.150 -24.580 70.410 -24.320 ;
        RECT 70.150 -24.930 70.410 -24.670 ;
        RECT 70.150 -28.190 70.410 -27.930 ;
        RECT 70.150 -28.540 70.410 -28.280 ;
        RECT 70.150 -31.800 70.410 -31.540 ;
        RECT 70.150 -32.150 70.410 -31.890 ;
        RECT 70.150 -35.410 70.410 -35.150 ;
        RECT 70.150 -35.760 70.410 -35.500 ;
        RECT 70.150 -39.020 70.410 -38.760 ;
        RECT 70.150 -39.370 70.410 -39.110 ;
        RECT 73.010 15.140 73.270 15.400 ;
        RECT 73.010 14.770 73.270 15.030 ;
        RECT 73.010 11.530 73.270 11.790 ;
        RECT 73.010 11.160 73.270 11.420 ;
        RECT 73.010 7.920 73.270 8.180 ;
        RECT 73.010 7.550 73.270 7.810 ;
        RECT 73.010 4.310 73.270 4.570 ;
        RECT 73.010 3.940 73.270 4.200 ;
        RECT 73.010 0.700 73.270 0.960 ;
        RECT 73.010 0.330 73.270 0.590 ;
        RECT 73.010 -2.910 73.270 -2.650 ;
        RECT 73.010 -3.280 73.270 -3.020 ;
        RECT 73.010 -6.520 73.270 -6.260 ;
        RECT 73.010 -6.890 73.270 -6.630 ;
        RECT 73.010 -10.130 73.270 -9.870 ;
        RECT 73.010 -10.500 73.270 -10.240 ;
        RECT 73.010 -13.740 73.270 -13.480 ;
        RECT 73.010 -14.110 73.270 -13.850 ;
        RECT 73.010 -17.350 73.270 -17.090 ;
        RECT 73.010 -17.720 73.270 -17.460 ;
        RECT 73.010 -20.960 73.270 -20.700 ;
        RECT 73.010 -21.330 73.270 -21.070 ;
        RECT 73.010 -24.570 73.270 -24.310 ;
        RECT 73.010 -24.940 73.270 -24.680 ;
        RECT 73.010 -28.180 73.270 -27.920 ;
        RECT 73.010 -28.550 73.270 -28.290 ;
        RECT 73.010 -31.790 73.270 -31.530 ;
        RECT 73.010 -32.160 73.270 -31.900 ;
        RECT 73.010 -35.400 73.270 -35.140 ;
        RECT 73.010 -35.770 73.270 -35.510 ;
        RECT 73.010 -39.010 73.270 -38.750 ;
        RECT 73.010 -39.380 73.270 -39.120 ;
        RECT 76.860 15.140 77.120 15.400 ;
        RECT 76.860 14.770 77.120 15.030 ;
        RECT 76.860 11.530 77.120 11.790 ;
        RECT 76.860 11.160 77.120 11.420 ;
        RECT 76.860 7.920 77.120 8.180 ;
        RECT 76.860 7.550 77.120 7.810 ;
        RECT 76.860 4.310 77.120 4.570 ;
        RECT 76.860 3.940 77.120 4.200 ;
        RECT 76.860 0.700 77.120 0.960 ;
        RECT 76.860 0.330 77.120 0.590 ;
        RECT 76.860 -2.910 77.120 -2.650 ;
        RECT 76.860 -3.280 77.120 -3.020 ;
        RECT 76.860 -6.520 77.120 -6.260 ;
        RECT 76.860 -6.890 77.120 -6.630 ;
        RECT 76.860 -10.130 77.120 -9.870 ;
        RECT 76.860 -10.500 77.120 -10.240 ;
        RECT 76.860 -13.740 77.120 -13.480 ;
        RECT 76.860 -14.110 77.120 -13.850 ;
        RECT 76.860 -17.350 77.120 -17.090 ;
        RECT 76.860 -17.720 77.120 -17.460 ;
        RECT 76.860 -20.960 77.120 -20.700 ;
        RECT 76.860 -21.330 77.120 -21.070 ;
        RECT 76.860 -24.570 77.120 -24.310 ;
        RECT 76.860 -24.940 77.120 -24.680 ;
        RECT 76.860 -28.180 77.120 -27.920 ;
        RECT 76.860 -28.550 77.120 -28.290 ;
        RECT 76.860 -31.790 77.120 -31.530 ;
        RECT 76.860 -32.160 77.120 -31.900 ;
        RECT 76.860 -35.400 77.120 -35.140 ;
        RECT 76.860 -35.770 77.120 -35.510 ;
        RECT 76.860 -39.010 77.120 -38.750 ;
        RECT 76.860 -39.380 77.120 -39.120 ;
        RECT 79.720 15.130 79.980 15.390 ;
        RECT 79.720 14.780 79.980 15.040 ;
        RECT 79.720 11.520 79.980 11.780 ;
        RECT 79.720 11.170 79.980 11.430 ;
        RECT 79.720 7.910 79.980 8.170 ;
        RECT 79.720 7.560 79.980 7.820 ;
        RECT 79.720 4.300 79.980 4.560 ;
        RECT 79.720 3.950 79.980 4.210 ;
        RECT 79.720 0.690 79.980 0.950 ;
        RECT 79.720 0.340 79.980 0.600 ;
        RECT 79.720 -2.920 79.980 -2.660 ;
        RECT 79.720 -3.270 79.980 -3.010 ;
        RECT 79.720 -6.530 79.980 -6.270 ;
        RECT 79.720 -6.880 79.980 -6.620 ;
        RECT 79.720 -10.140 79.980 -9.880 ;
        RECT 79.720 -10.490 79.980 -10.230 ;
        RECT 79.720 -13.750 79.980 -13.490 ;
        RECT 79.720 -14.100 79.980 -13.840 ;
        RECT 79.720 -17.360 79.980 -17.100 ;
        RECT 79.720 -17.710 79.980 -17.450 ;
        RECT 79.720 -20.970 79.980 -20.710 ;
        RECT 79.720 -21.320 79.980 -21.060 ;
        RECT 79.720 -24.580 79.980 -24.320 ;
        RECT 79.720 -24.930 79.980 -24.670 ;
        RECT 79.720 -28.190 79.980 -27.930 ;
        RECT 79.720 -28.540 79.980 -28.280 ;
        RECT 79.720 -31.800 79.980 -31.540 ;
        RECT 79.720 -32.150 79.980 -31.890 ;
        RECT 79.720 -35.410 79.980 -35.150 ;
        RECT 79.720 -35.760 79.980 -35.500 ;
        RECT 79.720 -39.020 79.980 -38.760 ;
        RECT 79.720 -39.370 79.980 -39.110 ;
        RECT 83.650 15.130 83.910 15.390 ;
        RECT 83.650 14.780 83.910 15.040 ;
        RECT 83.650 11.520 83.910 11.780 ;
        RECT 83.650 11.170 83.910 11.430 ;
        RECT 83.650 7.910 83.910 8.170 ;
        RECT 83.650 7.560 83.910 7.820 ;
        RECT 83.650 4.300 83.910 4.560 ;
        RECT 83.650 3.950 83.910 4.210 ;
        RECT 83.650 0.690 83.910 0.950 ;
        RECT 83.650 0.340 83.910 0.600 ;
        RECT 83.650 -2.920 83.910 -2.660 ;
        RECT 83.650 -3.270 83.910 -3.010 ;
        RECT 83.650 -6.530 83.910 -6.270 ;
        RECT 83.650 -6.880 83.910 -6.620 ;
        RECT 83.650 -10.140 83.910 -9.880 ;
        RECT 83.650 -10.490 83.910 -10.230 ;
        RECT 83.650 -13.750 83.910 -13.490 ;
        RECT 83.650 -14.100 83.910 -13.840 ;
        RECT 83.650 -17.360 83.910 -17.100 ;
        RECT 83.650 -17.710 83.910 -17.450 ;
        RECT 83.650 -20.970 83.910 -20.710 ;
        RECT 83.650 -21.320 83.910 -21.060 ;
        RECT 83.650 -24.580 83.910 -24.320 ;
        RECT 83.650 -24.930 83.910 -24.670 ;
        RECT 83.650 -28.190 83.910 -27.930 ;
        RECT 83.650 -28.540 83.910 -28.280 ;
        RECT 83.650 -31.800 83.910 -31.540 ;
        RECT 83.650 -32.150 83.910 -31.890 ;
        RECT 83.650 -35.410 83.910 -35.150 ;
        RECT 83.650 -35.760 83.910 -35.500 ;
        RECT 83.650 -39.020 83.910 -38.760 ;
        RECT 83.650 -39.370 83.910 -39.110 ;
        RECT 86.510 15.140 86.770 15.400 ;
        RECT 86.510 14.770 86.770 15.030 ;
        RECT 86.510 11.530 86.770 11.790 ;
        RECT 86.510 11.160 86.770 11.420 ;
        RECT 86.510 7.920 86.770 8.180 ;
        RECT 86.510 7.550 86.770 7.810 ;
        RECT 86.510 4.310 86.770 4.570 ;
        RECT 86.510 3.940 86.770 4.200 ;
        RECT 86.510 0.700 86.770 0.960 ;
        RECT 86.510 0.330 86.770 0.590 ;
        RECT 86.510 -2.910 86.770 -2.650 ;
        RECT 86.510 -3.280 86.770 -3.020 ;
        RECT 86.510 -6.520 86.770 -6.260 ;
        RECT 86.510 -6.890 86.770 -6.630 ;
        RECT 86.510 -10.130 86.770 -9.870 ;
        RECT 86.510 -10.500 86.770 -10.240 ;
        RECT 86.510 -13.740 86.770 -13.480 ;
        RECT 86.510 -14.110 86.770 -13.850 ;
        RECT 86.510 -17.350 86.770 -17.090 ;
        RECT 86.510 -17.720 86.770 -17.460 ;
        RECT 86.510 -20.960 86.770 -20.700 ;
        RECT 86.510 -21.330 86.770 -21.070 ;
        RECT 86.510 -24.570 86.770 -24.310 ;
        RECT 86.510 -24.940 86.770 -24.680 ;
        RECT 86.510 -28.180 86.770 -27.920 ;
        RECT 86.510 -28.550 86.770 -28.290 ;
        RECT 86.510 -31.790 86.770 -31.530 ;
        RECT 86.510 -32.160 86.770 -31.900 ;
        RECT 86.510 -35.400 86.770 -35.140 ;
        RECT 86.510 -35.770 86.770 -35.510 ;
        RECT 86.510 -39.010 86.770 -38.750 ;
        RECT 86.510 -39.380 86.770 -39.120 ;
        RECT 90.360 15.140 90.620 15.400 ;
        RECT 90.360 14.770 90.620 15.030 ;
        RECT 90.360 11.530 90.620 11.790 ;
        RECT 90.360 11.160 90.620 11.420 ;
        RECT 90.360 7.920 90.620 8.180 ;
        RECT 90.360 7.550 90.620 7.810 ;
        RECT 90.360 4.310 90.620 4.570 ;
        RECT 90.360 3.940 90.620 4.200 ;
        RECT 90.360 0.700 90.620 0.960 ;
        RECT 90.360 0.330 90.620 0.590 ;
        RECT 90.360 -2.910 90.620 -2.650 ;
        RECT 90.360 -3.280 90.620 -3.020 ;
        RECT 90.360 -6.520 90.620 -6.260 ;
        RECT 90.360 -6.890 90.620 -6.630 ;
        RECT 90.360 -10.130 90.620 -9.870 ;
        RECT 90.360 -10.500 90.620 -10.240 ;
        RECT 90.360 -13.740 90.620 -13.480 ;
        RECT 90.360 -14.110 90.620 -13.850 ;
        RECT 90.360 -17.350 90.620 -17.090 ;
        RECT 90.360 -17.720 90.620 -17.460 ;
        RECT 90.360 -20.960 90.620 -20.700 ;
        RECT 90.360 -21.330 90.620 -21.070 ;
        RECT 90.360 -24.570 90.620 -24.310 ;
        RECT 90.360 -24.940 90.620 -24.680 ;
        RECT 90.360 -28.180 90.620 -27.920 ;
        RECT 90.360 -28.550 90.620 -28.290 ;
        RECT 90.360 -31.790 90.620 -31.530 ;
        RECT 90.360 -32.160 90.620 -31.900 ;
        RECT 90.360 -35.400 90.620 -35.140 ;
        RECT 90.360 -35.770 90.620 -35.510 ;
        RECT 90.360 -39.010 90.620 -38.750 ;
        RECT 90.360 -39.380 90.620 -39.120 ;
        RECT 93.220 15.130 93.480 15.390 ;
        RECT 93.220 14.780 93.480 15.040 ;
        RECT 93.220 11.520 93.480 11.780 ;
        RECT 93.220 11.170 93.480 11.430 ;
        RECT 93.220 7.910 93.480 8.170 ;
        RECT 93.220 7.560 93.480 7.820 ;
        RECT 93.220 4.300 93.480 4.560 ;
        RECT 93.220 3.950 93.480 4.210 ;
        RECT 93.220 0.690 93.480 0.950 ;
        RECT 93.220 0.340 93.480 0.600 ;
        RECT 93.220 -2.920 93.480 -2.660 ;
        RECT 93.220 -3.270 93.480 -3.010 ;
        RECT 93.220 -6.530 93.480 -6.270 ;
        RECT 93.220 -6.880 93.480 -6.620 ;
        RECT 93.220 -10.140 93.480 -9.880 ;
        RECT 93.220 -10.490 93.480 -10.230 ;
        RECT 93.220 -13.750 93.480 -13.490 ;
        RECT 93.220 -14.100 93.480 -13.840 ;
        RECT 93.220 -17.360 93.480 -17.100 ;
        RECT 93.220 -17.710 93.480 -17.450 ;
        RECT 93.220 -20.970 93.480 -20.710 ;
        RECT 93.220 -21.320 93.480 -21.060 ;
        RECT 93.220 -24.580 93.480 -24.320 ;
        RECT 93.220 -24.930 93.480 -24.670 ;
        RECT 93.220 -28.190 93.480 -27.930 ;
        RECT 93.220 -28.540 93.480 -28.280 ;
        RECT 93.220 -31.800 93.480 -31.540 ;
        RECT 93.220 -32.150 93.480 -31.890 ;
        RECT 93.220 -35.410 93.480 -35.150 ;
        RECT 93.220 -35.760 93.480 -35.500 ;
        RECT 93.220 -39.020 93.480 -38.760 ;
        RECT 93.220 -39.370 93.480 -39.110 ;
        RECT 97.150 15.130 97.410 15.390 ;
        RECT 97.150 14.780 97.410 15.040 ;
        RECT 97.150 11.520 97.410 11.780 ;
        RECT 97.150 11.170 97.410 11.430 ;
        RECT 97.150 7.910 97.410 8.170 ;
        RECT 97.150 7.560 97.410 7.820 ;
        RECT 97.150 4.300 97.410 4.560 ;
        RECT 97.150 3.950 97.410 4.210 ;
        RECT 97.150 0.690 97.410 0.950 ;
        RECT 97.150 0.340 97.410 0.600 ;
        RECT 97.150 -2.920 97.410 -2.660 ;
        RECT 97.150 -3.270 97.410 -3.010 ;
        RECT 97.150 -6.530 97.410 -6.270 ;
        RECT 97.150 -6.880 97.410 -6.620 ;
        RECT 97.150 -10.140 97.410 -9.880 ;
        RECT 97.150 -10.490 97.410 -10.230 ;
        RECT 97.150 -13.750 97.410 -13.490 ;
        RECT 97.150 -14.100 97.410 -13.840 ;
        RECT 97.150 -17.360 97.410 -17.100 ;
        RECT 97.150 -17.710 97.410 -17.450 ;
        RECT 97.150 -20.970 97.410 -20.710 ;
        RECT 97.150 -21.320 97.410 -21.060 ;
        RECT 97.150 -24.580 97.410 -24.320 ;
        RECT 97.150 -24.930 97.410 -24.670 ;
        RECT 97.150 -28.190 97.410 -27.930 ;
        RECT 97.150 -28.540 97.410 -28.280 ;
        RECT 97.150 -31.800 97.410 -31.540 ;
        RECT 97.150 -32.150 97.410 -31.890 ;
        RECT 97.150 -35.410 97.410 -35.150 ;
        RECT 97.150 -35.760 97.410 -35.500 ;
        RECT 97.150 -39.020 97.410 -38.760 ;
        RECT 97.150 -39.370 97.410 -39.110 ;
        RECT 100.010 15.140 100.270 15.400 ;
        RECT 100.010 14.770 100.270 15.030 ;
        RECT 100.010 11.530 100.270 11.790 ;
        RECT 100.010 11.160 100.270 11.420 ;
        RECT 100.010 7.920 100.270 8.180 ;
        RECT 100.010 7.550 100.270 7.810 ;
        RECT 100.010 4.310 100.270 4.570 ;
        RECT 100.010 3.940 100.270 4.200 ;
        RECT 100.010 0.700 100.270 0.960 ;
        RECT 100.010 0.330 100.270 0.590 ;
        RECT 100.010 -2.910 100.270 -2.650 ;
        RECT 100.010 -3.280 100.270 -3.020 ;
        RECT 100.010 -6.520 100.270 -6.260 ;
        RECT 100.010 -6.890 100.270 -6.630 ;
        RECT 100.010 -10.130 100.270 -9.870 ;
        RECT 100.010 -10.500 100.270 -10.240 ;
        RECT 100.010 -13.740 100.270 -13.480 ;
        RECT 100.010 -14.110 100.270 -13.850 ;
        RECT 100.010 -17.350 100.270 -17.090 ;
        RECT 100.010 -17.720 100.270 -17.460 ;
        RECT 100.010 -20.960 100.270 -20.700 ;
        RECT 100.010 -21.330 100.270 -21.070 ;
        RECT 100.010 -24.570 100.270 -24.310 ;
        RECT 100.010 -24.940 100.270 -24.680 ;
        RECT 100.010 -28.180 100.270 -27.920 ;
        RECT 100.010 -28.550 100.270 -28.290 ;
        RECT 100.010 -31.790 100.270 -31.530 ;
        RECT 100.010 -32.160 100.270 -31.900 ;
        RECT 100.010 -35.400 100.270 -35.140 ;
        RECT 100.010 -35.770 100.270 -35.510 ;
        RECT 100.010 -39.010 100.270 -38.750 ;
        RECT 100.010 -39.380 100.270 -39.120 ;
        RECT 103.860 15.140 104.120 15.400 ;
        RECT 103.860 14.770 104.120 15.030 ;
        RECT 103.860 11.530 104.120 11.790 ;
        RECT 103.860 11.160 104.120 11.420 ;
        RECT 103.860 7.920 104.120 8.180 ;
        RECT 103.860 7.550 104.120 7.810 ;
        RECT 103.860 4.310 104.120 4.570 ;
        RECT 103.860 3.940 104.120 4.200 ;
        RECT 103.860 0.700 104.120 0.960 ;
        RECT 103.860 0.330 104.120 0.590 ;
        RECT 103.860 -2.910 104.120 -2.650 ;
        RECT 103.860 -3.280 104.120 -3.020 ;
        RECT 103.860 -6.520 104.120 -6.260 ;
        RECT 103.860 -6.890 104.120 -6.630 ;
        RECT 103.860 -10.130 104.120 -9.870 ;
        RECT 103.860 -10.500 104.120 -10.240 ;
        RECT 103.860 -13.740 104.120 -13.480 ;
        RECT 103.860 -14.110 104.120 -13.850 ;
        RECT 103.860 -17.350 104.120 -17.090 ;
        RECT 103.860 -17.720 104.120 -17.460 ;
        RECT 103.860 -20.960 104.120 -20.700 ;
        RECT 103.860 -21.330 104.120 -21.070 ;
        RECT 103.860 -24.570 104.120 -24.310 ;
        RECT 103.860 -24.940 104.120 -24.680 ;
        RECT 103.860 -28.180 104.120 -27.920 ;
        RECT 103.860 -28.550 104.120 -28.290 ;
        RECT 103.860 -31.790 104.120 -31.530 ;
        RECT 103.860 -32.160 104.120 -31.900 ;
        RECT 103.860 -35.400 104.120 -35.140 ;
        RECT 103.860 -35.770 104.120 -35.510 ;
        RECT 103.860 -39.010 104.120 -38.750 ;
        RECT 103.860 -39.380 104.120 -39.120 ;
        RECT 106.720 15.130 106.980 15.390 ;
        RECT 106.720 14.780 106.980 15.040 ;
        RECT 106.720 11.520 106.980 11.780 ;
        RECT 106.720 11.170 106.980 11.430 ;
        RECT 106.720 7.910 106.980 8.170 ;
        RECT 106.720 7.560 106.980 7.820 ;
        RECT 106.720 4.300 106.980 4.560 ;
        RECT 106.720 3.950 106.980 4.210 ;
        RECT 106.720 0.690 106.980 0.950 ;
        RECT 106.720 0.340 106.980 0.600 ;
        RECT 106.720 -2.920 106.980 -2.660 ;
        RECT 106.720 -3.270 106.980 -3.010 ;
        RECT 106.720 -6.530 106.980 -6.270 ;
        RECT 106.720 -6.880 106.980 -6.620 ;
        RECT 106.720 -10.140 106.980 -9.880 ;
        RECT 106.720 -10.490 106.980 -10.230 ;
        RECT 106.720 -13.750 106.980 -13.490 ;
        RECT 106.720 -14.100 106.980 -13.840 ;
        RECT 106.720 -17.360 106.980 -17.100 ;
        RECT 106.720 -17.710 106.980 -17.450 ;
        RECT 106.720 -20.970 106.980 -20.710 ;
        RECT 106.720 -21.320 106.980 -21.060 ;
        RECT 106.720 -24.580 106.980 -24.320 ;
        RECT 106.720 -24.930 106.980 -24.670 ;
        RECT 106.720 -28.190 106.980 -27.930 ;
        RECT 106.720 -28.540 106.980 -28.280 ;
        RECT 106.720 -31.800 106.980 -31.540 ;
        RECT 106.720 -32.150 106.980 -31.890 ;
        RECT 106.720 -35.410 106.980 -35.150 ;
        RECT 106.720 -35.760 106.980 -35.500 ;
        RECT 106.720 -39.020 106.980 -38.760 ;
        RECT 106.720 -39.370 106.980 -39.110 ;
        RECT 110.650 15.130 110.910 15.390 ;
        RECT 110.650 14.780 110.910 15.040 ;
        RECT 110.650 11.520 110.910 11.780 ;
        RECT 110.650 11.170 110.910 11.430 ;
        RECT 110.650 7.910 110.910 8.170 ;
        RECT 110.650 7.560 110.910 7.820 ;
        RECT 110.650 4.300 110.910 4.560 ;
        RECT 110.650 3.950 110.910 4.210 ;
        RECT 110.650 0.690 110.910 0.950 ;
        RECT 110.650 0.340 110.910 0.600 ;
        RECT 110.650 -2.920 110.910 -2.660 ;
        RECT 110.650 -3.270 110.910 -3.010 ;
        RECT 110.650 -6.530 110.910 -6.270 ;
        RECT 110.650 -6.880 110.910 -6.620 ;
        RECT 110.650 -10.140 110.910 -9.880 ;
        RECT 110.650 -10.490 110.910 -10.230 ;
        RECT 110.650 -13.750 110.910 -13.490 ;
        RECT 110.650 -14.100 110.910 -13.840 ;
        RECT 110.650 -17.360 110.910 -17.100 ;
        RECT 110.650 -17.710 110.910 -17.450 ;
        RECT 110.650 -20.970 110.910 -20.710 ;
        RECT 110.650 -21.320 110.910 -21.060 ;
        RECT 110.650 -24.580 110.910 -24.320 ;
        RECT 110.650 -24.930 110.910 -24.670 ;
        RECT 110.650 -28.190 110.910 -27.930 ;
        RECT 110.650 -28.540 110.910 -28.280 ;
        RECT 110.650 -31.800 110.910 -31.540 ;
        RECT 110.650 -32.150 110.910 -31.890 ;
        RECT 110.650 -35.410 110.910 -35.150 ;
        RECT 110.650 -35.760 110.910 -35.500 ;
        RECT 110.650 -39.020 110.910 -38.760 ;
        RECT 110.650 -39.370 110.910 -39.110 ;
        RECT 113.510 15.140 113.770 15.400 ;
        RECT 113.510 14.770 113.770 15.030 ;
        RECT 113.510 11.530 113.770 11.790 ;
        RECT 113.510 11.160 113.770 11.420 ;
        RECT 113.510 7.920 113.770 8.180 ;
        RECT 113.510 7.550 113.770 7.810 ;
        RECT 113.510 4.310 113.770 4.570 ;
        RECT 113.510 3.940 113.770 4.200 ;
        RECT 113.510 0.700 113.770 0.960 ;
        RECT 113.510 0.330 113.770 0.590 ;
        RECT 113.510 -2.910 113.770 -2.650 ;
        RECT 113.510 -3.280 113.770 -3.020 ;
        RECT 113.510 -6.520 113.770 -6.260 ;
        RECT 113.510 -6.890 113.770 -6.630 ;
        RECT 113.510 -10.130 113.770 -9.870 ;
        RECT 113.510 -10.500 113.770 -10.240 ;
        RECT 113.510 -13.740 113.770 -13.480 ;
        RECT 113.510 -14.110 113.770 -13.850 ;
        RECT 113.510 -17.350 113.770 -17.090 ;
        RECT 113.510 -17.720 113.770 -17.460 ;
        RECT 113.510 -20.960 113.770 -20.700 ;
        RECT 113.510 -21.330 113.770 -21.070 ;
        RECT 113.510 -24.570 113.770 -24.310 ;
        RECT 113.510 -24.940 113.770 -24.680 ;
        RECT 113.510 -28.180 113.770 -27.920 ;
        RECT 113.510 -28.550 113.770 -28.290 ;
        RECT 113.510 -31.790 113.770 -31.530 ;
        RECT 113.510 -32.160 113.770 -31.900 ;
        RECT 113.510 -35.400 113.770 -35.140 ;
        RECT 113.510 -35.770 113.770 -35.510 ;
        RECT 113.510 -39.010 113.770 -38.750 ;
        RECT 113.510 -39.380 113.770 -39.120 ;
        RECT 117.360 15.140 117.620 15.400 ;
        RECT 117.360 14.770 117.620 15.030 ;
        RECT 117.360 11.530 117.620 11.790 ;
        RECT 117.360 11.160 117.620 11.420 ;
        RECT 117.360 7.920 117.620 8.180 ;
        RECT 117.360 7.550 117.620 7.810 ;
        RECT 117.360 4.310 117.620 4.570 ;
        RECT 117.360 3.940 117.620 4.200 ;
        RECT 117.360 0.700 117.620 0.960 ;
        RECT 117.360 0.330 117.620 0.590 ;
        RECT 117.360 -2.910 117.620 -2.650 ;
        RECT 117.360 -3.280 117.620 -3.020 ;
        RECT 117.360 -6.520 117.620 -6.260 ;
        RECT 117.360 -6.890 117.620 -6.630 ;
        RECT 117.360 -10.130 117.620 -9.870 ;
        RECT 117.360 -10.500 117.620 -10.240 ;
        RECT 117.360 -13.740 117.620 -13.480 ;
        RECT 117.360 -14.110 117.620 -13.850 ;
        RECT 117.360 -17.350 117.620 -17.090 ;
        RECT 117.360 -17.720 117.620 -17.460 ;
        RECT 117.360 -20.960 117.620 -20.700 ;
        RECT 117.360 -21.330 117.620 -21.070 ;
        RECT 117.360 -24.570 117.620 -24.310 ;
        RECT 117.360 -24.940 117.620 -24.680 ;
        RECT 117.360 -28.180 117.620 -27.920 ;
        RECT 117.360 -28.550 117.620 -28.290 ;
        RECT 117.360 -31.790 117.620 -31.530 ;
        RECT 117.360 -32.160 117.620 -31.900 ;
        RECT 117.360 -35.400 117.620 -35.140 ;
        RECT 117.360 -35.770 117.620 -35.510 ;
        RECT 117.360 -39.010 117.620 -38.750 ;
        RECT 117.360 -39.380 117.620 -39.120 ;
        RECT 120.220 15.130 120.480 15.390 ;
        RECT 120.220 14.780 120.480 15.040 ;
        RECT 120.220 11.520 120.480 11.780 ;
        RECT 120.220 11.170 120.480 11.430 ;
        RECT 120.220 7.910 120.480 8.170 ;
        RECT 120.220 7.560 120.480 7.820 ;
        RECT 120.220 4.300 120.480 4.560 ;
        RECT 120.220 3.950 120.480 4.210 ;
        RECT 120.220 0.690 120.480 0.950 ;
        RECT 120.220 0.340 120.480 0.600 ;
        RECT 120.220 -2.920 120.480 -2.660 ;
        RECT 120.220 -3.270 120.480 -3.010 ;
        RECT 120.220 -6.530 120.480 -6.270 ;
        RECT 120.220 -6.880 120.480 -6.620 ;
        RECT 120.220 -10.140 120.480 -9.880 ;
        RECT 120.220 -10.490 120.480 -10.230 ;
        RECT 120.220 -13.750 120.480 -13.490 ;
        RECT 120.220 -14.100 120.480 -13.840 ;
        RECT 120.220 -17.360 120.480 -17.100 ;
        RECT 120.220 -17.710 120.480 -17.450 ;
        RECT 120.220 -20.970 120.480 -20.710 ;
        RECT 120.220 -21.320 120.480 -21.060 ;
        RECT 120.220 -24.580 120.480 -24.320 ;
        RECT 120.220 -24.930 120.480 -24.670 ;
        RECT 120.220 -28.190 120.480 -27.930 ;
        RECT 120.220 -28.540 120.480 -28.280 ;
        RECT 120.220 -31.800 120.480 -31.540 ;
        RECT 120.220 -32.150 120.480 -31.890 ;
        RECT 120.220 -35.410 120.480 -35.150 ;
        RECT 120.220 -35.760 120.480 -35.500 ;
        RECT 120.220 -39.020 120.480 -38.760 ;
        RECT 120.220 -39.370 120.480 -39.110 ;
        RECT 124.150 15.130 124.410 15.390 ;
        RECT 124.150 14.780 124.410 15.040 ;
        RECT 124.150 11.520 124.410 11.780 ;
        RECT 124.150 11.170 124.410 11.430 ;
        RECT 124.150 7.910 124.410 8.170 ;
        RECT 124.150 7.560 124.410 7.820 ;
        RECT 124.150 4.300 124.410 4.560 ;
        RECT 124.150 3.950 124.410 4.210 ;
        RECT 124.150 0.690 124.410 0.950 ;
        RECT 124.150 0.340 124.410 0.600 ;
        RECT 124.150 -2.920 124.410 -2.660 ;
        RECT 124.150 -3.270 124.410 -3.010 ;
        RECT 124.150 -6.530 124.410 -6.270 ;
        RECT 124.150 -6.880 124.410 -6.620 ;
        RECT 124.150 -10.140 124.410 -9.880 ;
        RECT 124.150 -10.490 124.410 -10.230 ;
        RECT 124.150 -13.750 124.410 -13.490 ;
        RECT 124.150 -14.100 124.410 -13.840 ;
        RECT 124.150 -17.360 124.410 -17.100 ;
        RECT 124.150 -17.710 124.410 -17.450 ;
        RECT 124.150 -20.970 124.410 -20.710 ;
        RECT 124.150 -21.320 124.410 -21.060 ;
        RECT 124.150 -24.580 124.410 -24.320 ;
        RECT 124.150 -24.930 124.410 -24.670 ;
        RECT 124.150 -28.190 124.410 -27.930 ;
        RECT 124.150 -28.540 124.410 -28.280 ;
        RECT 124.150 -31.800 124.410 -31.540 ;
        RECT 124.150 -32.150 124.410 -31.890 ;
        RECT 124.150 -35.410 124.410 -35.150 ;
        RECT 124.150 -35.760 124.410 -35.500 ;
        RECT 124.150 -39.020 124.410 -38.760 ;
        RECT 124.150 -39.370 124.410 -39.110 ;
        RECT 127.010 15.140 127.270 15.400 ;
        RECT 127.010 14.770 127.270 15.030 ;
        RECT 127.010 11.530 127.270 11.790 ;
        RECT 127.010 11.160 127.270 11.420 ;
        RECT 127.010 7.920 127.270 8.180 ;
        RECT 127.010 7.550 127.270 7.810 ;
        RECT 127.010 4.310 127.270 4.570 ;
        RECT 127.010 3.940 127.270 4.200 ;
        RECT 127.010 0.700 127.270 0.960 ;
        RECT 127.010 0.330 127.270 0.590 ;
        RECT 127.010 -2.910 127.270 -2.650 ;
        RECT 127.010 -3.280 127.270 -3.020 ;
        RECT 127.010 -6.520 127.270 -6.260 ;
        RECT 127.010 -6.890 127.270 -6.630 ;
        RECT 127.010 -10.130 127.270 -9.870 ;
        RECT 127.010 -10.500 127.270 -10.240 ;
        RECT 127.010 -13.740 127.270 -13.480 ;
        RECT 127.010 -14.110 127.270 -13.850 ;
        RECT 127.010 -17.350 127.270 -17.090 ;
        RECT 127.010 -17.720 127.270 -17.460 ;
        RECT 127.010 -20.960 127.270 -20.700 ;
        RECT 127.010 -21.330 127.270 -21.070 ;
        RECT 127.010 -24.570 127.270 -24.310 ;
        RECT 127.010 -24.940 127.270 -24.680 ;
        RECT 127.010 -28.180 127.270 -27.920 ;
        RECT 127.010 -28.550 127.270 -28.290 ;
        RECT 127.010 -31.790 127.270 -31.530 ;
        RECT 127.010 -32.160 127.270 -31.900 ;
        RECT 127.010 -35.400 127.270 -35.140 ;
        RECT 127.010 -35.770 127.270 -35.510 ;
        RECT 127.010 -39.010 127.270 -38.750 ;
        RECT 127.010 -39.380 127.270 -39.120 ;
        RECT 130.860 15.140 131.120 15.400 ;
        RECT 130.860 14.770 131.120 15.030 ;
        RECT 130.860 11.530 131.120 11.790 ;
        RECT 130.860 11.160 131.120 11.420 ;
        RECT 130.860 7.920 131.120 8.180 ;
        RECT 130.860 7.550 131.120 7.810 ;
        RECT 130.860 4.310 131.120 4.570 ;
        RECT 130.860 3.940 131.120 4.200 ;
        RECT 130.860 0.700 131.120 0.960 ;
        RECT 130.860 0.330 131.120 0.590 ;
        RECT 130.860 -2.910 131.120 -2.650 ;
        RECT 130.860 -3.280 131.120 -3.020 ;
        RECT 130.860 -6.520 131.120 -6.260 ;
        RECT 130.860 -6.890 131.120 -6.630 ;
        RECT 130.860 -10.130 131.120 -9.870 ;
        RECT 130.860 -10.500 131.120 -10.240 ;
        RECT 130.860 -13.740 131.120 -13.480 ;
        RECT 130.860 -14.110 131.120 -13.850 ;
        RECT 130.860 -17.350 131.120 -17.090 ;
        RECT 130.860 -17.720 131.120 -17.460 ;
        RECT 130.860 -20.960 131.120 -20.700 ;
        RECT 130.860 -21.330 131.120 -21.070 ;
        RECT 130.860 -24.570 131.120 -24.310 ;
        RECT 130.860 -24.940 131.120 -24.680 ;
        RECT 130.860 -28.180 131.120 -27.920 ;
        RECT 130.860 -28.550 131.120 -28.290 ;
        RECT 130.860 -31.790 131.120 -31.530 ;
        RECT 130.860 -32.160 131.120 -31.900 ;
        RECT 130.860 -35.400 131.120 -35.140 ;
        RECT 130.860 -35.770 131.120 -35.510 ;
        RECT 130.860 -39.010 131.120 -38.750 ;
        RECT 130.860 -39.380 131.120 -39.120 ;
        RECT 133.720 15.130 133.980 15.390 ;
        RECT 133.720 14.780 133.980 15.040 ;
        RECT 133.720 11.520 133.980 11.780 ;
        RECT 133.720 11.170 133.980 11.430 ;
        RECT 133.720 7.910 133.980 8.170 ;
        RECT 133.720 7.560 133.980 7.820 ;
        RECT 133.720 4.300 133.980 4.560 ;
        RECT 133.720 3.950 133.980 4.210 ;
        RECT 133.720 0.690 133.980 0.950 ;
        RECT 133.720 0.340 133.980 0.600 ;
        RECT 133.720 -2.920 133.980 -2.660 ;
        RECT 133.720 -3.270 133.980 -3.010 ;
        RECT 133.720 -6.530 133.980 -6.270 ;
        RECT 133.720 -6.880 133.980 -6.620 ;
        RECT 133.720 -10.140 133.980 -9.880 ;
        RECT 133.720 -10.490 133.980 -10.230 ;
        RECT 133.720 -13.750 133.980 -13.490 ;
        RECT 133.720 -14.100 133.980 -13.840 ;
        RECT 133.720 -17.360 133.980 -17.100 ;
        RECT 133.720 -17.710 133.980 -17.450 ;
        RECT 133.720 -20.970 133.980 -20.710 ;
        RECT 133.720 -21.320 133.980 -21.060 ;
        RECT 133.720 -24.580 133.980 -24.320 ;
        RECT 133.720 -24.930 133.980 -24.670 ;
        RECT 133.720 -28.190 133.980 -27.930 ;
        RECT 133.720 -28.540 133.980 -28.280 ;
        RECT 133.720 -31.800 133.980 -31.540 ;
        RECT 133.720 -32.150 133.980 -31.890 ;
        RECT 133.720 -35.410 133.980 -35.150 ;
        RECT 133.720 -35.760 133.980 -35.500 ;
        RECT 133.720 -39.020 133.980 -38.760 ;
        RECT 133.720 -39.370 133.980 -39.110 ;
        RECT 137.650 15.130 137.910 15.390 ;
        RECT 137.650 14.780 137.910 15.040 ;
        RECT 137.650 11.520 137.910 11.780 ;
        RECT 137.650 11.170 137.910 11.430 ;
        RECT 137.650 7.910 137.910 8.170 ;
        RECT 137.650 7.560 137.910 7.820 ;
        RECT 137.650 4.300 137.910 4.560 ;
        RECT 137.650 3.950 137.910 4.210 ;
        RECT 137.650 0.690 137.910 0.950 ;
        RECT 137.650 0.340 137.910 0.600 ;
        RECT 137.650 -2.920 137.910 -2.660 ;
        RECT 137.650 -3.270 137.910 -3.010 ;
        RECT 137.650 -6.530 137.910 -6.270 ;
        RECT 137.650 -6.880 137.910 -6.620 ;
        RECT 137.650 -10.140 137.910 -9.880 ;
        RECT 137.650 -10.490 137.910 -10.230 ;
        RECT 137.650 -13.750 137.910 -13.490 ;
        RECT 137.650 -14.100 137.910 -13.840 ;
        RECT 137.650 -17.360 137.910 -17.100 ;
        RECT 137.650 -17.710 137.910 -17.450 ;
        RECT 137.650 -20.970 137.910 -20.710 ;
        RECT 137.650 -21.320 137.910 -21.060 ;
        RECT 137.650 -24.580 137.910 -24.320 ;
        RECT 137.650 -24.930 137.910 -24.670 ;
        RECT 137.650 -28.190 137.910 -27.930 ;
        RECT 137.650 -28.540 137.910 -28.280 ;
        RECT 137.650 -31.800 137.910 -31.540 ;
        RECT 137.650 -32.150 137.910 -31.890 ;
        RECT 137.650 -35.410 137.910 -35.150 ;
        RECT 137.650 -35.760 137.910 -35.500 ;
        RECT 137.650 -39.020 137.910 -38.760 ;
        RECT 137.650 -39.370 137.910 -39.110 ;
        RECT 140.510 15.140 140.770 15.400 ;
        RECT 140.510 14.770 140.770 15.030 ;
        RECT 140.510 11.530 140.770 11.790 ;
        RECT 140.510 11.160 140.770 11.420 ;
        RECT 140.510 7.920 140.770 8.180 ;
        RECT 140.510 7.550 140.770 7.810 ;
        RECT 140.510 4.310 140.770 4.570 ;
        RECT 140.510 3.940 140.770 4.200 ;
        RECT 140.510 0.700 140.770 0.960 ;
        RECT 140.510 0.330 140.770 0.590 ;
        RECT 140.510 -2.910 140.770 -2.650 ;
        RECT 140.510 -3.280 140.770 -3.020 ;
        RECT 140.510 -6.520 140.770 -6.260 ;
        RECT 140.510 -6.890 140.770 -6.630 ;
        RECT 140.510 -10.130 140.770 -9.870 ;
        RECT 140.510 -10.500 140.770 -10.240 ;
        RECT 140.510 -13.740 140.770 -13.480 ;
        RECT 140.510 -14.110 140.770 -13.850 ;
        RECT 140.510 -17.350 140.770 -17.090 ;
        RECT 140.510 -17.720 140.770 -17.460 ;
        RECT 140.510 -20.960 140.770 -20.700 ;
        RECT 140.510 -21.330 140.770 -21.070 ;
        RECT 140.510 -24.570 140.770 -24.310 ;
        RECT 140.510 -24.940 140.770 -24.680 ;
        RECT 140.510 -28.180 140.770 -27.920 ;
        RECT 140.510 -28.550 140.770 -28.290 ;
        RECT 140.510 -31.790 140.770 -31.530 ;
        RECT 140.510 -32.160 140.770 -31.900 ;
        RECT 140.510 -35.400 140.770 -35.140 ;
        RECT 140.510 -35.770 140.770 -35.510 ;
        RECT 140.510 -39.010 140.770 -38.750 ;
        RECT 140.510 -39.380 140.770 -39.120 ;
        RECT 144.360 15.140 144.620 15.400 ;
        RECT 144.360 14.770 144.620 15.030 ;
        RECT 144.360 11.530 144.620 11.790 ;
        RECT 144.360 11.160 144.620 11.420 ;
        RECT 144.360 7.920 144.620 8.180 ;
        RECT 144.360 7.550 144.620 7.810 ;
        RECT 144.360 4.310 144.620 4.570 ;
        RECT 144.360 3.940 144.620 4.200 ;
        RECT 144.360 0.700 144.620 0.960 ;
        RECT 144.360 0.330 144.620 0.590 ;
        RECT 144.360 -2.910 144.620 -2.650 ;
        RECT 144.360 -3.280 144.620 -3.020 ;
        RECT 144.360 -6.520 144.620 -6.260 ;
        RECT 144.360 -6.890 144.620 -6.630 ;
        RECT 144.360 -10.130 144.620 -9.870 ;
        RECT 144.360 -10.500 144.620 -10.240 ;
        RECT 144.360 -13.740 144.620 -13.480 ;
        RECT 144.360 -14.110 144.620 -13.850 ;
        RECT 144.360 -17.350 144.620 -17.090 ;
        RECT 144.360 -17.720 144.620 -17.460 ;
        RECT 144.360 -20.960 144.620 -20.700 ;
        RECT 144.360 -21.330 144.620 -21.070 ;
        RECT 144.360 -24.570 144.620 -24.310 ;
        RECT 144.360 -24.940 144.620 -24.680 ;
        RECT 144.360 -28.180 144.620 -27.920 ;
        RECT 144.360 -28.550 144.620 -28.290 ;
        RECT 144.360 -31.790 144.620 -31.530 ;
        RECT 144.360 -32.160 144.620 -31.900 ;
        RECT 144.360 -35.400 144.620 -35.140 ;
        RECT 144.360 -35.770 144.620 -35.510 ;
        RECT 144.360 -39.010 144.620 -38.750 ;
        RECT 144.360 -39.380 144.620 -39.120 ;
        RECT 147.220 15.130 147.480 15.390 ;
        RECT 147.220 14.780 147.480 15.040 ;
        RECT 147.220 11.520 147.480 11.780 ;
        RECT 147.220 11.170 147.480 11.430 ;
        RECT 147.220 7.910 147.480 8.170 ;
        RECT 147.220 7.560 147.480 7.820 ;
        RECT 147.220 4.300 147.480 4.560 ;
        RECT 147.220 3.950 147.480 4.210 ;
        RECT 147.220 0.690 147.480 0.950 ;
        RECT 147.220 0.340 147.480 0.600 ;
        RECT 147.220 -2.920 147.480 -2.660 ;
        RECT 147.220 -3.270 147.480 -3.010 ;
        RECT 147.220 -6.530 147.480 -6.270 ;
        RECT 147.220 -6.880 147.480 -6.620 ;
        RECT 147.220 -10.140 147.480 -9.880 ;
        RECT 147.220 -10.490 147.480 -10.230 ;
        RECT 147.220 -13.750 147.480 -13.490 ;
        RECT 147.220 -14.100 147.480 -13.840 ;
        RECT 147.220 -17.360 147.480 -17.100 ;
        RECT 147.220 -17.710 147.480 -17.450 ;
        RECT 147.220 -20.970 147.480 -20.710 ;
        RECT 147.220 -21.320 147.480 -21.060 ;
        RECT 147.220 -24.580 147.480 -24.320 ;
        RECT 147.220 -24.930 147.480 -24.670 ;
        RECT 147.220 -28.190 147.480 -27.930 ;
        RECT 147.220 -28.540 147.480 -28.280 ;
        RECT 147.220 -31.800 147.480 -31.540 ;
        RECT 147.220 -32.150 147.480 -31.890 ;
        RECT 147.220 -35.410 147.480 -35.150 ;
        RECT 147.220 -35.760 147.480 -35.500 ;
        RECT 147.220 -39.020 147.480 -38.760 ;
        RECT 147.220 -39.370 147.480 -39.110 ;
        RECT 151.150 15.130 151.410 15.390 ;
        RECT 151.150 14.780 151.410 15.040 ;
        RECT 151.150 11.520 151.410 11.780 ;
        RECT 151.150 11.170 151.410 11.430 ;
        RECT 151.150 7.910 151.410 8.170 ;
        RECT 151.150 7.560 151.410 7.820 ;
        RECT 151.150 4.300 151.410 4.560 ;
        RECT 151.150 3.950 151.410 4.210 ;
        RECT 151.150 0.690 151.410 0.950 ;
        RECT 151.150 0.340 151.410 0.600 ;
        RECT 151.150 -2.920 151.410 -2.660 ;
        RECT 151.150 -3.270 151.410 -3.010 ;
        RECT 151.150 -6.530 151.410 -6.270 ;
        RECT 151.150 -6.880 151.410 -6.620 ;
        RECT 151.150 -10.140 151.410 -9.880 ;
        RECT 151.150 -10.490 151.410 -10.230 ;
        RECT 151.150 -13.750 151.410 -13.490 ;
        RECT 151.150 -14.100 151.410 -13.840 ;
        RECT 151.150 -17.360 151.410 -17.100 ;
        RECT 151.150 -17.710 151.410 -17.450 ;
        RECT 151.150 -20.970 151.410 -20.710 ;
        RECT 151.150 -21.320 151.410 -21.060 ;
        RECT 151.150 -24.580 151.410 -24.320 ;
        RECT 151.150 -24.930 151.410 -24.670 ;
        RECT 151.150 -28.190 151.410 -27.930 ;
        RECT 151.150 -28.540 151.410 -28.280 ;
        RECT 151.150 -31.800 151.410 -31.540 ;
        RECT 151.150 -32.150 151.410 -31.890 ;
        RECT 151.150 -35.410 151.410 -35.150 ;
        RECT 151.150 -35.760 151.410 -35.500 ;
        RECT 151.150 -39.020 151.410 -38.760 ;
        RECT 151.150 -39.370 151.410 -39.110 ;
        RECT 154.010 15.140 154.270 15.400 ;
        RECT 154.010 14.770 154.270 15.030 ;
        RECT 154.010 11.530 154.270 11.790 ;
        RECT 154.010 11.160 154.270 11.420 ;
        RECT 154.010 7.920 154.270 8.180 ;
        RECT 154.010 7.550 154.270 7.810 ;
        RECT 154.010 4.310 154.270 4.570 ;
        RECT 154.010 3.940 154.270 4.200 ;
        RECT 154.010 0.700 154.270 0.960 ;
        RECT 154.010 0.330 154.270 0.590 ;
        RECT 154.010 -2.910 154.270 -2.650 ;
        RECT 154.010 -3.280 154.270 -3.020 ;
        RECT 154.010 -6.520 154.270 -6.260 ;
        RECT 154.010 -6.890 154.270 -6.630 ;
        RECT 154.010 -10.130 154.270 -9.870 ;
        RECT 154.010 -10.500 154.270 -10.240 ;
        RECT 154.010 -13.740 154.270 -13.480 ;
        RECT 154.010 -14.110 154.270 -13.850 ;
        RECT 154.010 -17.350 154.270 -17.090 ;
        RECT 154.010 -17.720 154.270 -17.460 ;
        RECT 154.010 -20.960 154.270 -20.700 ;
        RECT 154.010 -21.330 154.270 -21.070 ;
        RECT 154.010 -24.570 154.270 -24.310 ;
        RECT 154.010 -24.940 154.270 -24.680 ;
        RECT 154.010 -28.180 154.270 -27.920 ;
        RECT 154.010 -28.550 154.270 -28.290 ;
        RECT 154.010 -31.790 154.270 -31.530 ;
        RECT 154.010 -32.160 154.270 -31.900 ;
        RECT 154.010 -35.400 154.270 -35.140 ;
        RECT 154.010 -35.770 154.270 -35.510 ;
        RECT 154.010 -39.010 154.270 -38.750 ;
        RECT 154.010 -39.380 154.270 -39.120 ;
        RECT 157.860 15.140 158.120 15.400 ;
        RECT 157.860 14.770 158.120 15.030 ;
        RECT 157.860 11.530 158.120 11.790 ;
        RECT 157.860 11.160 158.120 11.420 ;
        RECT 157.860 7.920 158.120 8.180 ;
        RECT 157.860 7.550 158.120 7.810 ;
        RECT 157.860 4.310 158.120 4.570 ;
        RECT 157.860 3.940 158.120 4.200 ;
        RECT 157.860 0.700 158.120 0.960 ;
        RECT 157.860 0.330 158.120 0.590 ;
        RECT 157.860 -2.910 158.120 -2.650 ;
        RECT 157.860 -3.280 158.120 -3.020 ;
        RECT 157.860 -6.520 158.120 -6.260 ;
        RECT 157.860 -6.890 158.120 -6.630 ;
        RECT 157.860 -10.130 158.120 -9.870 ;
        RECT 157.860 -10.500 158.120 -10.240 ;
        RECT 157.860 -13.740 158.120 -13.480 ;
        RECT 157.860 -14.110 158.120 -13.850 ;
        RECT 157.860 -17.350 158.120 -17.090 ;
        RECT 157.860 -17.720 158.120 -17.460 ;
        RECT 157.860 -20.960 158.120 -20.700 ;
        RECT 157.860 -21.330 158.120 -21.070 ;
        RECT 157.860 -24.570 158.120 -24.310 ;
        RECT 157.860 -24.940 158.120 -24.680 ;
        RECT 157.860 -28.180 158.120 -27.920 ;
        RECT 157.860 -28.550 158.120 -28.290 ;
        RECT 157.860 -31.790 158.120 -31.530 ;
        RECT 157.860 -32.160 158.120 -31.900 ;
        RECT 157.860 -35.400 158.120 -35.140 ;
        RECT 157.860 -35.770 158.120 -35.510 ;
        RECT 157.860 -39.010 158.120 -38.750 ;
        RECT 157.860 -39.380 158.120 -39.120 ;
        RECT 160.720 15.130 160.980 15.390 ;
        RECT 160.720 14.780 160.980 15.040 ;
        RECT 160.720 11.520 160.980 11.780 ;
        RECT 160.720 11.170 160.980 11.430 ;
        RECT 160.720 7.910 160.980 8.170 ;
        RECT 160.720 7.560 160.980 7.820 ;
        RECT 160.720 4.300 160.980 4.560 ;
        RECT 160.720 3.950 160.980 4.210 ;
        RECT 160.720 0.690 160.980 0.950 ;
        RECT 160.720 0.340 160.980 0.600 ;
        RECT 160.720 -2.920 160.980 -2.660 ;
        RECT 160.720 -3.270 160.980 -3.010 ;
        RECT 160.720 -6.530 160.980 -6.270 ;
        RECT 160.720 -6.880 160.980 -6.620 ;
        RECT 160.720 -10.140 160.980 -9.880 ;
        RECT 160.720 -10.490 160.980 -10.230 ;
        RECT 160.720 -13.750 160.980 -13.490 ;
        RECT 160.720 -14.100 160.980 -13.840 ;
        RECT 160.720 -17.360 160.980 -17.100 ;
        RECT 160.720 -17.710 160.980 -17.450 ;
        RECT 160.720 -20.970 160.980 -20.710 ;
        RECT 160.720 -21.320 160.980 -21.060 ;
        RECT 160.720 -24.580 160.980 -24.320 ;
        RECT 160.720 -24.930 160.980 -24.670 ;
        RECT 160.720 -28.190 160.980 -27.930 ;
        RECT 160.720 -28.540 160.980 -28.280 ;
        RECT 160.720 -31.800 160.980 -31.540 ;
        RECT 160.720 -32.150 160.980 -31.890 ;
        RECT 160.720 -35.410 160.980 -35.150 ;
        RECT 160.720 -35.760 160.980 -35.500 ;
        RECT 160.720 -39.020 160.980 -38.760 ;
        RECT 160.720 -39.370 160.980 -39.110 ;
        RECT 164.650 15.130 164.910 15.390 ;
        RECT 164.650 14.780 164.910 15.040 ;
        RECT 164.650 11.520 164.910 11.780 ;
        RECT 164.650 11.170 164.910 11.430 ;
        RECT 164.650 7.910 164.910 8.170 ;
        RECT 164.650 7.560 164.910 7.820 ;
        RECT 164.650 4.300 164.910 4.560 ;
        RECT 164.650 3.950 164.910 4.210 ;
        RECT 164.650 0.690 164.910 0.950 ;
        RECT 164.650 0.340 164.910 0.600 ;
        RECT 164.650 -2.920 164.910 -2.660 ;
        RECT 164.650 -3.270 164.910 -3.010 ;
        RECT 164.650 -6.530 164.910 -6.270 ;
        RECT 164.650 -6.880 164.910 -6.620 ;
        RECT 164.650 -10.140 164.910 -9.880 ;
        RECT 164.650 -10.490 164.910 -10.230 ;
        RECT 164.650 -13.750 164.910 -13.490 ;
        RECT 164.650 -14.100 164.910 -13.840 ;
        RECT 164.650 -17.360 164.910 -17.100 ;
        RECT 164.650 -17.710 164.910 -17.450 ;
        RECT 164.650 -20.970 164.910 -20.710 ;
        RECT 164.650 -21.320 164.910 -21.060 ;
        RECT 164.650 -24.580 164.910 -24.320 ;
        RECT 164.650 -24.930 164.910 -24.670 ;
        RECT 164.650 -28.190 164.910 -27.930 ;
        RECT 164.650 -28.540 164.910 -28.280 ;
        RECT 164.650 -31.800 164.910 -31.540 ;
        RECT 164.650 -32.150 164.910 -31.890 ;
        RECT 164.650 -35.410 164.910 -35.150 ;
        RECT 164.650 -35.760 164.910 -35.500 ;
        RECT 164.650 -39.020 164.910 -38.760 ;
        RECT 164.650 -39.370 164.910 -39.110 ;
        RECT 167.510 15.140 167.770 15.400 ;
        RECT 167.510 14.770 167.770 15.030 ;
        RECT 167.510 11.530 167.770 11.790 ;
        RECT 167.510 11.160 167.770 11.420 ;
        RECT 167.510 7.920 167.770 8.180 ;
        RECT 167.510 7.550 167.770 7.810 ;
        RECT 167.510 4.310 167.770 4.570 ;
        RECT 167.510 3.940 167.770 4.200 ;
        RECT 167.510 0.700 167.770 0.960 ;
        RECT 167.510 0.330 167.770 0.590 ;
        RECT 167.510 -2.910 167.770 -2.650 ;
        RECT 167.510 -3.280 167.770 -3.020 ;
        RECT 167.510 -6.520 167.770 -6.260 ;
        RECT 167.510 -6.890 167.770 -6.630 ;
        RECT 167.510 -10.130 167.770 -9.870 ;
        RECT 167.510 -10.500 167.770 -10.240 ;
        RECT 167.510 -13.740 167.770 -13.480 ;
        RECT 167.510 -14.110 167.770 -13.850 ;
        RECT 167.510 -17.350 167.770 -17.090 ;
        RECT 167.510 -17.720 167.770 -17.460 ;
        RECT 167.510 -20.960 167.770 -20.700 ;
        RECT 167.510 -21.330 167.770 -21.070 ;
        RECT 167.510 -24.570 167.770 -24.310 ;
        RECT 167.510 -24.940 167.770 -24.680 ;
        RECT 167.510 -28.180 167.770 -27.920 ;
        RECT 167.510 -28.550 167.770 -28.290 ;
        RECT 167.510 -31.790 167.770 -31.530 ;
        RECT 167.510 -32.160 167.770 -31.900 ;
        RECT 167.510 -35.400 167.770 -35.140 ;
        RECT 167.510 -35.770 167.770 -35.510 ;
        RECT 167.510 -39.010 167.770 -38.750 ;
        RECT 167.510 -39.380 167.770 -39.120 ;
        RECT 171.360 15.140 171.620 15.400 ;
        RECT 171.360 14.770 171.620 15.030 ;
        RECT 171.360 11.530 171.620 11.790 ;
        RECT 171.360 11.160 171.620 11.420 ;
        RECT 171.360 7.920 171.620 8.180 ;
        RECT 171.360 7.550 171.620 7.810 ;
        RECT 171.360 4.310 171.620 4.570 ;
        RECT 171.360 3.940 171.620 4.200 ;
        RECT 171.360 0.700 171.620 0.960 ;
        RECT 171.360 0.330 171.620 0.590 ;
        RECT 171.360 -2.910 171.620 -2.650 ;
        RECT 171.360 -3.280 171.620 -3.020 ;
        RECT 171.360 -6.520 171.620 -6.260 ;
        RECT 171.360 -6.890 171.620 -6.630 ;
        RECT 171.360 -10.130 171.620 -9.870 ;
        RECT 171.360 -10.500 171.620 -10.240 ;
        RECT 171.360 -13.740 171.620 -13.480 ;
        RECT 171.360 -14.110 171.620 -13.850 ;
        RECT 171.360 -17.350 171.620 -17.090 ;
        RECT 171.360 -17.720 171.620 -17.460 ;
        RECT 171.360 -20.960 171.620 -20.700 ;
        RECT 171.360 -21.330 171.620 -21.070 ;
        RECT 171.360 -24.570 171.620 -24.310 ;
        RECT 171.360 -24.940 171.620 -24.680 ;
        RECT 171.360 -28.180 171.620 -27.920 ;
        RECT 171.360 -28.550 171.620 -28.290 ;
        RECT 171.360 -31.790 171.620 -31.530 ;
        RECT 171.360 -32.160 171.620 -31.900 ;
        RECT 171.360 -35.400 171.620 -35.140 ;
        RECT 171.360 -35.770 171.620 -35.510 ;
        RECT 171.360 -39.010 171.620 -38.750 ;
        RECT 171.360 -39.380 171.620 -39.120 ;
        RECT 174.220 15.130 174.480 15.390 ;
        RECT 174.220 14.780 174.480 15.040 ;
        RECT 174.220 11.520 174.480 11.780 ;
        RECT 174.220 11.170 174.480 11.430 ;
        RECT 174.220 7.910 174.480 8.170 ;
        RECT 174.220 7.560 174.480 7.820 ;
        RECT 174.220 4.300 174.480 4.560 ;
        RECT 174.220 3.950 174.480 4.210 ;
        RECT 174.220 0.690 174.480 0.950 ;
        RECT 174.220 0.340 174.480 0.600 ;
        RECT 174.220 -2.920 174.480 -2.660 ;
        RECT 174.220 -3.270 174.480 -3.010 ;
        RECT 174.220 -6.530 174.480 -6.270 ;
        RECT 174.220 -6.880 174.480 -6.620 ;
        RECT 174.220 -10.140 174.480 -9.880 ;
        RECT 174.220 -10.490 174.480 -10.230 ;
        RECT 174.220 -13.750 174.480 -13.490 ;
        RECT 174.220 -14.100 174.480 -13.840 ;
        RECT 174.220 -17.360 174.480 -17.100 ;
        RECT 174.220 -17.710 174.480 -17.450 ;
        RECT 174.220 -20.970 174.480 -20.710 ;
        RECT 174.220 -21.320 174.480 -21.060 ;
        RECT 174.220 -24.580 174.480 -24.320 ;
        RECT 174.220 -24.930 174.480 -24.670 ;
        RECT 174.220 -28.190 174.480 -27.930 ;
        RECT 174.220 -28.540 174.480 -28.280 ;
        RECT 174.220 -31.800 174.480 -31.540 ;
        RECT 174.220 -32.150 174.480 -31.890 ;
        RECT 174.220 -35.410 174.480 -35.150 ;
        RECT 174.220 -35.760 174.480 -35.500 ;
        RECT 174.220 -39.020 174.480 -38.760 ;
        RECT 174.220 -39.370 174.480 -39.110 ;
        RECT 178.150 15.130 178.410 15.390 ;
        RECT 178.150 14.780 178.410 15.040 ;
        RECT 178.150 11.520 178.410 11.780 ;
        RECT 178.150 11.170 178.410 11.430 ;
        RECT 178.150 7.910 178.410 8.170 ;
        RECT 178.150 7.560 178.410 7.820 ;
        RECT 178.150 4.300 178.410 4.560 ;
        RECT 178.150 3.950 178.410 4.210 ;
        RECT 178.150 0.690 178.410 0.950 ;
        RECT 178.150 0.340 178.410 0.600 ;
        RECT 178.150 -2.920 178.410 -2.660 ;
        RECT 178.150 -3.270 178.410 -3.010 ;
        RECT 178.150 -6.530 178.410 -6.270 ;
        RECT 178.150 -6.880 178.410 -6.620 ;
        RECT 178.150 -10.140 178.410 -9.880 ;
        RECT 178.150 -10.490 178.410 -10.230 ;
        RECT 178.150 -13.750 178.410 -13.490 ;
        RECT 178.150 -14.100 178.410 -13.840 ;
        RECT 178.150 -17.360 178.410 -17.100 ;
        RECT 178.150 -17.710 178.410 -17.450 ;
        RECT 178.150 -20.970 178.410 -20.710 ;
        RECT 178.150 -21.320 178.410 -21.060 ;
        RECT 178.150 -24.580 178.410 -24.320 ;
        RECT 178.150 -24.930 178.410 -24.670 ;
        RECT 178.150 -28.190 178.410 -27.930 ;
        RECT 178.150 -28.540 178.410 -28.280 ;
        RECT 178.150 -31.800 178.410 -31.540 ;
        RECT 178.150 -32.150 178.410 -31.890 ;
        RECT 178.150 -35.410 178.410 -35.150 ;
        RECT 178.150 -35.760 178.410 -35.500 ;
        RECT 178.150 -39.020 178.410 -38.760 ;
        RECT 178.150 -39.370 178.410 -39.110 ;
        RECT 181.010 15.140 181.270 15.400 ;
        RECT 181.010 14.770 181.270 15.030 ;
        RECT 181.010 11.530 181.270 11.790 ;
        RECT 181.010 11.160 181.270 11.420 ;
        RECT 181.010 7.920 181.270 8.180 ;
        RECT 181.010 7.550 181.270 7.810 ;
        RECT 181.010 4.310 181.270 4.570 ;
        RECT 181.010 3.940 181.270 4.200 ;
        RECT 181.010 0.700 181.270 0.960 ;
        RECT 181.010 0.330 181.270 0.590 ;
        RECT 181.010 -2.910 181.270 -2.650 ;
        RECT 181.010 -3.280 181.270 -3.020 ;
        RECT 181.010 -6.520 181.270 -6.260 ;
        RECT 181.010 -6.890 181.270 -6.630 ;
        RECT 181.010 -10.130 181.270 -9.870 ;
        RECT 181.010 -10.500 181.270 -10.240 ;
        RECT 181.010 -13.740 181.270 -13.480 ;
        RECT 181.010 -14.110 181.270 -13.850 ;
        RECT 181.010 -17.350 181.270 -17.090 ;
        RECT 181.010 -17.720 181.270 -17.460 ;
        RECT 181.010 -20.960 181.270 -20.700 ;
        RECT 181.010 -21.330 181.270 -21.070 ;
        RECT 181.010 -24.570 181.270 -24.310 ;
        RECT 181.010 -24.940 181.270 -24.680 ;
        RECT 181.010 -28.180 181.270 -27.920 ;
        RECT 181.010 -28.550 181.270 -28.290 ;
        RECT 181.010 -31.790 181.270 -31.530 ;
        RECT 181.010 -32.160 181.270 -31.900 ;
        RECT 181.010 -35.400 181.270 -35.140 ;
        RECT 181.010 -35.770 181.270 -35.510 ;
        RECT 181.010 -39.010 181.270 -38.750 ;
        RECT 181.010 -39.380 181.270 -39.120 ;
        RECT 184.860 15.140 185.120 15.400 ;
        RECT 184.860 14.770 185.120 15.030 ;
        RECT 184.860 11.530 185.120 11.790 ;
        RECT 184.860 11.160 185.120 11.420 ;
        RECT 184.860 7.920 185.120 8.180 ;
        RECT 184.860 7.550 185.120 7.810 ;
        RECT 184.860 4.310 185.120 4.570 ;
        RECT 184.860 3.940 185.120 4.200 ;
        RECT 184.860 0.700 185.120 0.960 ;
        RECT 184.860 0.330 185.120 0.590 ;
        RECT 184.860 -2.910 185.120 -2.650 ;
        RECT 184.860 -3.280 185.120 -3.020 ;
        RECT 184.860 -6.520 185.120 -6.260 ;
        RECT 184.860 -6.890 185.120 -6.630 ;
        RECT 184.860 -10.130 185.120 -9.870 ;
        RECT 184.860 -10.500 185.120 -10.240 ;
        RECT 184.860 -13.740 185.120 -13.480 ;
        RECT 184.860 -14.110 185.120 -13.850 ;
        RECT 184.860 -17.350 185.120 -17.090 ;
        RECT 184.860 -17.720 185.120 -17.460 ;
        RECT 184.860 -20.960 185.120 -20.700 ;
        RECT 184.860 -21.330 185.120 -21.070 ;
        RECT 184.860 -24.570 185.120 -24.310 ;
        RECT 184.860 -24.940 185.120 -24.680 ;
        RECT 184.860 -28.180 185.120 -27.920 ;
        RECT 184.860 -28.550 185.120 -28.290 ;
        RECT 184.860 -31.790 185.120 -31.530 ;
        RECT 184.860 -32.160 185.120 -31.900 ;
        RECT 184.860 -35.400 185.120 -35.140 ;
        RECT 184.860 -35.770 185.120 -35.510 ;
        RECT 184.860 -39.010 185.120 -38.750 ;
        RECT 184.860 -39.380 185.120 -39.120 ;
        RECT 187.720 15.130 187.980 15.390 ;
        RECT 187.720 14.780 187.980 15.040 ;
        RECT 187.720 11.520 187.980 11.780 ;
        RECT 187.720 11.170 187.980 11.430 ;
        RECT 187.720 7.910 187.980 8.170 ;
        RECT 187.720 7.560 187.980 7.820 ;
        RECT 187.720 4.300 187.980 4.560 ;
        RECT 187.720 3.950 187.980 4.210 ;
        RECT 187.720 0.690 187.980 0.950 ;
        RECT 187.720 0.340 187.980 0.600 ;
        RECT 187.720 -2.920 187.980 -2.660 ;
        RECT 187.720 -3.270 187.980 -3.010 ;
        RECT 187.720 -6.530 187.980 -6.270 ;
        RECT 187.720 -6.880 187.980 -6.620 ;
        RECT 187.720 -10.140 187.980 -9.880 ;
        RECT 187.720 -10.490 187.980 -10.230 ;
        RECT 187.720 -13.750 187.980 -13.490 ;
        RECT 187.720 -14.100 187.980 -13.840 ;
        RECT 187.720 -17.360 187.980 -17.100 ;
        RECT 187.720 -17.710 187.980 -17.450 ;
        RECT 187.720 -20.970 187.980 -20.710 ;
        RECT 187.720 -21.320 187.980 -21.060 ;
        RECT 187.720 -24.580 187.980 -24.320 ;
        RECT 187.720 -24.930 187.980 -24.670 ;
        RECT 187.720 -28.190 187.980 -27.930 ;
        RECT 187.720 -28.540 187.980 -28.280 ;
        RECT 187.720 -31.800 187.980 -31.540 ;
        RECT 187.720 -32.150 187.980 -31.890 ;
        RECT 187.720 -35.410 187.980 -35.150 ;
        RECT 187.720 -35.760 187.980 -35.500 ;
        RECT 187.720 -39.020 187.980 -38.760 ;
        RECT 187.720 -39.370 187.980 -39.110 ;
        RECT 191.650 15.130 191.910 15.390 ;
        RECT 191.650 14.780 191.910 15.040 ;
        RECT 191.650 11.520 191.910 11.780 ;
        RECT 191.650 11.170 191.910 11.430 ;
        RECT 191.650 7.910 191.910 8.170 ;
        RECT 191.650 7.560 191.910 7.820 ;
        RECT 191.650 4.300 191.910 4.560 ;
        RECT 191.650 3.950 191.910 4.210 ;
        RECT 191.650 0.690 191.910 0.950 ;
        RECT 191.650 0.340 191.910 0.600 ;
        RECT 191.650 -2.920 191.910 -2.660 ;
        RECT 191.650 -3.270 191.910 -3.010 ;
        RECT 191.650 -6.530 191.910 -6.270 ;
        RECT 191.650 -6.880 191.910 -6.620 ;
        RECT 191.650 -10.140 191.910 -9.880 ;
        RECT 191.650 -10.490 191.910 -10.230 ;
        RECT 191.650 -13.750 191.910 -13.490 ;
        RECT 191.650 -14.100 191.910 -13.840 ;
        RECT 191.650 -17.360 191.910 -17.100 ;
        RECT 191.650 -17.710 191.910 -17.450 ;
        RECT 191.650 -20.970 191.910 -20.710 ;
        RECT 191.650 -21.320 191.910 -21.060 ;
        RECT 191.650 -24.580 191.910 -24.320 ;
        RECT 191.650 -24.930 191.910 -24.670 ;
        RECT 191.650 -28.190 191.910 -27.930 ;
        RECT 191.650 -28.540 191.910 -28.280 ;
        RECT 191.650 -31.800 191.910 -31.540 ;
        RECT 191.650 -32.150 191.910 -31.890 ;
        RECT 191.650 -35.410 191.910 -35.150 ;
        RECT 191.650 -35.760 191.910 -35.500 ;
        RECT 191.650 -39.020 191.910 -38.760 ;
        RECT 191.650 -39.370 191.910 -39.110 ;
        RECT 194.510 15.140 194.770 15.400 ;
        RECT 194.510 14.770 194.770 15.030 ;
        RECT 194.510 11.530 194.770 11.790 ;
        RECT 194.510 11.160 194.770 11.420 ;
        RECT 194.510 7.920 194.770 8.180 ;
        RECT 194.510 7.550 194.770 7.810 ;
        RECT 194.510 4.310 194.770 4.570 ;
        RECT 194.510 3.940 194.770 4.200 ;
        RECT 194.510 0.700 194.770 0.960 ;
        RECT 194.510 0.330 194.770 0.590 ;
        RECT 194.510 -2.910 194.770 -2.650 ;
        RECT 194.510 -3.280 194.770 -3.020 ;
        RECT 194.510 -6.520 194.770 -6.260 ;
        RECT 194.510 -6.890 194.770 -6.630 ;
        RECT 194.510 -10.130 194.770 -9.870 ;
        RECT 194.510 -10.500 194.770 -10.240 ;
        RECT 194.510 -13.740 194.770 -13.480 ;
        RECT 194.510 -14.110 194.770 -13.850 ;
        RECT 194.510 -17.350 194.770 -17.090 ;
        RECT 194.510 -17.720 194.770 -17.460 ;
        RECT 194.510 -20.960 194.770 -20.700 ;
        RECT 194.510 -21.330 194.770 -21.070 ;
        RECT 194.510 -24.570 194.770 -24.310 ;
        RECT 194.510 -24.940 194.770 -24.680 ;
        RECT 194.510 -28.180 194.770 -27.920 ;
        RECT 194.510 -28.550 194.770 -28.290 ;
        RECT 194.510 -31.790 194.770 -31.530 ;
        RECT 194.510 -32.160 194.770 -31.900 ;
        RECT 194.510 -35.400 194.770 -35.140 ;
        RECT 194.510 -35.770 194.770 -35.510 ;
        RECT 194.510 -39.010 194.770 -38.750 ;
        RECT 194.510 -39.380 194.770 -39.120 ;
        RECT 198.360 15.140 198.620 15.400 ;
        RECT 198.360 14.770 198.620 15.030 ;
        RECT 198.360 11.530 198.620 11.790 ;
        RECT 198.360 11.160 198.620 11.420 ;
        RECT 198.360 7.920 198.620 8.180 ;
        RECT 198.360 7.550 198.620 7.810 ;
        RECT 198.360 4.310 198.620 4.570 ;
        RECT 198.360 3.940 198.620 4.200 ;
        RECT 198.360 0.700 198.620 0.960 ;
        RECT 198.360 0.330 198.620 0.590 ;
        RECT 198.360 -2.910 198.620 -2.650 ;
        RECT 198.360 -3.280 198.620 -3.020 ;
        RECT 198.360 -6.520 198.620 -6.260 ;
        RECT 198.360 -6.890 198.620 -6.630 ;
        RECT 198.360 -10.130 198.620 -9.870 ;
        RECT 198.360 -10.500 198.620 -10.240 ;
        RECT 198.360 -13.740 198.620 -13.480 ;
        RECT 198.360 -14.110 198.620 -13.850 ;
        RECT 198.360 -17.350 198.620 -17.090 ;
        RECT 198.360 -17.720 198.620 -17.460 ;
        RECT 198.360 -20.960 198.620 -20.700 ;
        RECT 198.360 -21.330 198.620 -21.070 ;
        RECT 198.360 -24.570 198.620 -24.310 ;
        RECT 198.360 -24.940 198.620 -24.680 ;
        RECT 198.360 -28.180 198.620 -27.920 ;
        RECT 198.360 -28.550 198.620 -28.290 ;
        RECT 198.360 -31.790 198.620 -31.530 ;
        RECT 198.360 -32.160 198.620 -31.900 ;
        RECT 198.360 -35.400 198.620 -35.140 ;
        RECT 198.360 -35.770 198.620 -35.510 ;
        RECT 198.360 -39.010 198.620 -38.750 ;
        RECT 198.360 -39.380 198.620 -39.120 ;
        RECT 201.220 15.130 201.480 15.390 ;
        RECT 201.220 14.780 201.480 15.040 ;
        RECT 201.220 11.520 201.480 11.780 ;
        RECT 201.220 11.170 201.480 11.430 ;
        RECT 201.220 7.910 201.480 8.170 ;
        RECT 201.220 7.560 201.480 7.820 ;
        RECT 201.220 4.300 201.480 4.560 ;
        RECT 201.220 3.950 201.480 4.210 ;
        RECT 201.220 0.690 201.480 0.950 ;
        RECT 201.220 0.340 201.480 0.600 ;
        RECT 201.220 -2.920 201.480 -2.660 ;
        RECT 201.220 -3.270 201.480 -3.010 ;
        RECT 201.220 -6.530 201.480 -6.270 ;
        RECT 201.220 -6.880 201.480 -6.620 ;
        RECT 201.220 -10.140 201.480 -9.880 ;
        RECT 201.220 -10.490 201.480 -10.230 ;
        RECT 201.220 -13.750 201.480 -13.490 ;
        RECT 201.220 -14.100 201.480 -13.840 ;
        RECT 201.220 -17.360 201.480 -17.100 ;
        RECT 201.220 -17.710 201.480 -17.450 ;
        RECT 201.220 -20.970 201.480 -20.710 ;
        RECT 201.220 -21.320 201.480 -21.060 ;
        RECT 201.220 -24.580 201.480 -24.320 ;
        RECT 201.220 -24.930 201.480 -24.670 ;
        RECT 201.220 -28.190 201.480 -27.930 ;
        RECT 201.220 -28.540 201.480 -28.280 ;
        RECT 201.220 -31.800 201.480 -31.540 ;
        RECT 201.220 -32.150 201.480 -31.890 ;
        RECT 201.220 -35.410 201.480 -35.150 ;
        RECT 201.220 -35.760 201.480 -35.500 ;
        RECT 201.220 -39.020 201.480 -38.760 ;
        RECT 201.220 -39.370 201.480 -39.110 ;
        RECT 205.150 15.130 205.410 15.390 ;
        RECT 205.150 14.780 205.410 15.040 ;
        RECT 205.150 11.520 205.410 11.780 ;
        RECT 205.150 11.170 205.410 11.430 ;
        RECT 205.150 7.910 205.410 8.170 ;
        RECT 205.150 7.560 205.410 7.820 ;
        RECT 205.150 4.300 205.410 4.560 ;
        RECT 205.150 3.950 205.410 4.210 ;
        RECT 205.150 0.690 205.410 0.950 ;
        RECT 205.150 0.340 205.410 0.600 ;
        RECT 205.150 -2.920 205.410 -2.660 ;
        RECT 205.150 -3.270 205.410 -3.010 ;
        RECT 205.150 -6.530 205.410 -6.270 ;
        RECT 205.150 -6.880 205.410 -6.620 ;
        RECT 205.150 -10.140 205.410 -9.880 ;
        RECT 205.150 -10.490 205.410 -10.230 ;
        RECT 205.150 -13.750 205.410 -13.490 ;
        RECT 205.150 -14.100 205.410 -13.840 ;
        RECT 205.150 -17.360 205.410 -17.100 ;
        RECT 205.150 -17.710 205.410 -17.450 ;
        RECT 205.150 -20.970 205.410 -20.710 ;
        RECT 205.150 -21.320 205.410 -21.060 ;
        RECT 205.150 -24.580 205.410 -24.320 ;
        RECT 205.150 -24.930 205.410 -24.670 ;
        RECT 205.150 -28.190 205.410 -27.930 ;
        RECT 205.150 -28.540 205.410 -28.280 ;
        RECT 205.150 -31.800 205.410 -31.540 ;
        RECT 205.150 -32.150 205.410 -31.890 ;
        RECT 205.150 -35.410 205.410 -35.150 ;
        RECT 205.150 -35.760 205.410 -35.500 ;
        RECT 205.150 -39.020 205.410 -38.760 ;
        RECT 205.150 -39.370 205.410 -39.110 ;
        RECT 208.010 15.140 208.270 15.400 ;
        RECT 208.010 14.770 208.270 15.030 ;
        RECT 208.010 11.530 208.270 11.790 ;
        RECT 208.010 11.160 208.270 11.420 ;
        RECT 208.010 7.920 208.270 8.180 ;
        RECT 208.010 7.550 208.270 7.810 ;
        RECT 208.010 4.310 208.270 4.570 ;
        RECT 208.010 3.940 208.270 4.200 ;
        RECT 208.010 0.700 208.270 0.960 ;
        RECT 208.010 0.330 208.270 0.590 ;
        RECT 208.010 -2.910 208.270 -2.650 ;
        RECT 208.010 -3.280 208.270 -3.020 ;
        RECT 208.010 -6.520 208.270 -6.260 ;
        RECT 208.010 -6.890 208.270 -6.630 ;
        RECT 208.010 -10.130 208.270 -9.870 ;
        RECT 208.010 -10.500 208.270 -10.240 ;
        RECT 208.010 -13.740 208.270 -13.480 ;
        RECT 208.010 -14.110 208.270 -13.850 ;
        RECT 208.010 -17.350 208.270 -17.090 ;
        RECT 208.010 -17.720 208.270 -17.460 ;
        RECT 208.010 -20.960 208.270 -20.700 ;
        RECT 208.010 -21.330 208.270 -21.070 ;
        RECT 208.010 -24.570 208.270 -24.310 ;
        RECT 208.010 -24.940 208.270 -24.680 ;
        RECT 208.010 -28.180 208.270 -27.920 ;
        RECT 208.010 -28.550 208.270 -28.290 ;
        RECT 208.010 -31.790 208.270 -31.530 ;
        RECT 208.010 -32.160 208.270 -31.900 ;
        RECT 208.010 -35.400 208.270 -35.140 ;
        RECT 208.010 -35.770 208.270 -35.510 ;
        RECT 208.010 -39.010 208.270 -38.750 ;
        RECT 208.010 -39.380 208.270 -39.120 ;
        RECT 211.860 15.140 212.120 15.400 ;
        RECT 211.860 14.770 212.120 15.030 ;
        RECT 211.860 11.530 212.120 11.790 ;
        RECT 211.860 11.160 212.120 11.420 ;
        RECT 211.860 7.920 212.120 8.180 ;
        RECT 211.860 7.550 212.120 7.810 ;
        RECT 211.860 4.310 212.120 4.570 ;
        RECT 211.860 3.940 212.120 4.200 ;
        RECT 211.860 0.700 212.120 0.960 ;
        RECT 211.860 0.330 212.120 0.590 ;
        RECT 211.860 -2.910 212.120 -2.650 ;
        RECT 211.860 -3.280 212.120 -3.020 ;
        RECT 211.860 -6.520 212.120 -6.260 ;
        RECT 211.860 -6.890 212.120 -6.630 ;
        RECT 211.860 -10.130 212.120 -9.870 ;
        RECT 211.860 -10.500 212.120 -10.240 ;
        RECT 211.860 -13.740 212.120 -13.480 ;
        RECT 211.860 -14.110 212.120 -13.850 ;
        RECT 211.860 -17.350 212.120 -17.090 ;
        RECT 211.860 -17.720 212.120 -17.460 ;
        RECT 211.860 -20.960 212.120 -20.700 ;
        RECT 211.860 -21.330 212.120 -21.070 ;
        RECT 211.860 -24.570 212.120 -24.310 ;
        RECT 211.860 -24.940 212.120 -24.680 ;
        RECT 211.860 -28.180 212.120 -27.920 ;
        RECT 211.860 -28.550 212.120 -28.290 ;
        RECT 211.860 -31.790 212.120 -31.530 ;
        RECT 211.860 -32.160 212.120 -31.900 ;
        RECT 211.860 -35.400 212.120 -35.140 ;
        RECT 211.860 -35.770 212.120 -35.510 ;
        RECT 211.860 -39.010 212.120 -38.750 ;
        RECT 211.860 -39.380 212.120 -39.120 ;
        RECT 214.720 15.130 214.980 15.390 ;
        RECT 214.720 14.780 214.980 15.040 ;
        RECT 214.720 11.520 214.980 11.780 ;
        RECT 214.720 11.170 214.980 11.430 ;
        RECT 214.720 7.910 214.980 8.170 ;
        RECT 214.720 7.560 214.980 7.820 ;
        RECT 214.720 4.300 214.980 4.560 ;
        RECT 214.720 3.950 214.980 4.210 ;
        RECT 214.720 0.690 214.980 0.950 ;
        RECT 214.720 0.340 214.980 0.600 ;
        RECT 214.720 -2.920 214.980 -2.660 ;
        RECT 214.720 -3.270 214.980 -3.010 ;
        RECT 214.720 -6.530 214.980 -6.270 ;
        RECT 214.720 -6.880 214.980 -6.620 ;
        RECT 214.720 -10.140 214.980 -9.880 ;
        RECT 214.720 -10.490 214.980 -10.230 ;
        RECT 214.720 -13.750 214.980 -13.490 ;
        RECT 214.720 -14.100 214.980 -13.840 ;
        RECT 214.720 -17.360 214.980 -17.100 ;
        RECT 214.720 -17.710 214.980 -17.450 ;
        RECT 214.720 -20.970 214.980 -20.710 ;
        RECT 214.720 -21.320 214.980 -21.060 ;
        RECT 214.720 -24.580 214.980 -24.320 ;
        RECT 214.720 -24.930 214.980 -24.670 ;
        RECT 214.720 -28.190 214.980 -27.930 ;
        RECT 214.720 -28.540 214.980 -28.280 ;
        RECT 214.720 -31.800 214.980 -31.540 ;
        RECT 214.720 -32.150 214.980 -31.890 ;
        RECT 214.720 -35.410 214.980 -35.150 ;
        RECT 214.720 -35.760 214.980 -35.500 ;
        RECT 214.720 -39.020 214.980 -38.760 ;
        RECT 214.720 -39.370 214.980 -39.110 ;
      LAYER met2 ;
        RECT 9.260 15.410 9.710 15.500 ;
        RECT 12.110 15.410 12.570 15.490 ;
        RECT 9.260 15.180 12.570 15.410 ;
        RECT 9.260 14.990 9.710 15.180 ;
        RECT 12.110 14.990 12.570 15.180 ;
        RECT 9.260 14.760 12.570 14.990 ;
        RECT 9.260 14.670 9.710 14.760 ;
        RECT 12.110 14.680 12.570 14.760 ;
        RECT 16.060 15.410 16.520 15.490 ;
        RECT 18.920 15.410 19.370 15.500 ;
        RECT 16.060 15.180 19.370 15.410 ;
        RECT 16.060 14.990 16.520 15.180 ;
        RECT 18.920 14.990 19.370 15.180 ;
        RECT 16.060 14.760 19.370 14.990 ;
        RECT 16.060 14.680 16.520 14.760 ;
        RECT 18.920 14.670 19.370 14.760 ;
        RECT 22.760 15.410 23.210 15.500 ;
        RECT 25.610 15.410 26.070 15.490 ;
        RECT 22.760 15.180 26.070 15.410 ;
        RECT 22.760 14.990 23.210 15.180 ;
        RECT 25.610 14.990 26.070 15.180 ;
        RECT 22.760 14.760 26.070 14.990 ;
        RECT 22.760 14.670 23.210 14.760 ;
        RECT 25.610 14.680 26.070 14.760 ;
        RECT 29.560 15.410 30.020 15.490 ;
        RECT 32.420 15.410 32.870 15.500 ;
        RECT 29.560 15.180 32.870 15.410 ;
        RECT 29.560 14.990 30.020 15.180 ;
        RECT 32.420 14.990 32.870 15.180 ;
        RECT 29.560 14.760 32.870 14.990 ;
        RECT 29.560 14.680 30.020 14.760 ;
        RECT 32.420 14.670 32.870 14.760 ;
        RECT 36.260 15.410 36.710 15.500 ;
        RECT 39.110 15.410 39.570 15.490 ;
        RECT 36.260 15.180 39.570 15.410 ;
        RECT 36.260 14.990 36.710 15.180 ;
        RECT 39.110 14.990 39.570 15.180 ;
        RECT 36.260 14.760 39.570 14.990 ;
        RECT 36.260 14.670 36.710 14.760 ;
        RECT 39.110 14.680 39.570 14.760 ;
        RECT 43.060 15.410 43.520 15.490 ;
        RECT 45.920 15.410 46.370 15.500 ;
        RECT 43.060 15.180 46.370 15.410 ;
        RECT 43.060 14.990 43.520 15.180 ;
        RECT 45.920 14.990 46.370 15.180 ;
        RECT 43.060 14.760 46.370 14.990 ;
        RECT 43.060 14.680 43.520 14.760 ;
        RECT 45.920 14.670 46.370 14.760 ;
        RECT 49.760 15.410 50.210 15.500 ;
        RECT 52.610 15.410 53.070 15.490 ;
        RECT 49.760 15.180 53.070 15.410 ;
        RECT 49.760 14.990 50.210 15.180 ;
        RECT 52.610 14.990 53.070 15.180 ;
        RECT 49.760 14.760 53.070 14.990 ;
        RECT 49.760 14.670 50.210 14.760 ;
        RECT 52.610 14.680 53.070 14.760 ;
        RECT 56.560 15.410 57.020 15.490 ;
        RECT 59.420 15.410 59.870 15.500 ;
        RECT 56.560 15.180 59.870 15.410 ;
        RECT 56.560 14.990 57.020 15.180 ;
        RECT 59.420 14.990 59.870 15.180 ;
        RECT 56.560 14.760 59.870 14.990 ;
        RECT 56.560 14.680 57.020 14.760 ;
        RECT 59.420 14.670 59.870 14.760 ;
        RECT 63.260 15.410 63.710 15.500 ;
        RECT 66.110 15.410 66.570 15.490 ;
        RECT 63.260 15.180 66.570 15.410 ;
        RECT 63.260 14.990 63.710 15.180 ;
        RECT 66.110 14.990 66.570 15.180 ;
        RECT 63.260 14.760 66.570 14.990 ;
        RECT 63.260 14.670 63.710 14.760 ;
        RECT 66.110 14.680 66.570 14.760 ;
        RECT 70.060 15.410 70.520 15.490 ;
        RECT 72.920 15.410 73.370 15.500 ;
        RECT 70.060 15.180 73.370 15.410 ;
        RECT 70.060 14.990 70.520 15.180 ;
        RECT 72.920 14.990 73.370 15.180 ;
        RECT 70.060 14.760 73.370 14.990 ;
        RECT 70.060 14.680 70.520 14.760 ;
        RECT 72.920 14.670 73.370 14.760 ;
        RECT 76.760 15.410 77.210 15.500 ;
        RECT 79.610 15.410 80.070 15.490 ;
        RECT 76.760 15.180 80.070 15.410 ;
        RECT 76.760 14.990 77.210 15.180 ;
        RECT 79.610 14.990 80.070 15.180 ;
        RECT 76.760 14.760 80.070 14.990 ;
        RECT 76.760 14.670 77.210 14.760 ;
        RECT 79.610 14.680 80.070 14.760 ;
        RECT 83.560 15.410 84.020 15.490 ;
        RECT 86.420 15.410 86.870 15.500 ;
        RECT 83.560 15.180 86.870 15.410 ;
        RECT 83.560 14.990 84.020 15.180 ;
        RECT 86.420 14.990 86.870 15.180 ;
        RECT 83.560 14.760 86.870 14.990 ;
        RECT 83.560 14.680 84.020 14.760 ;
        RECT 86.420 14.670 86.870 14.760 ;
        RECT 90.260 15.410 90.710 15.500 ;
        RECT 93.110 15.410 93.570 15.490 ;
        RECT 90.260 15.180 93.570 15.410 ;
        RECT 90.260 14.990 90.710 15.180 ;
        RECT 93.110 14.990 93.570 15.180 ;
        RECT 90.260 14.760 93.570 14.990 ;
        RECT 90.260 14.670 90.710 14.760 ;
        RECT 93.110 14.680 93.570 14.760 ;
        RECT 97.060 15.410 97.520 15.490 ;
        RECT 99.920 15.410 100.370 15.500 ;
        RECT 97.060 15.180 100.370 15.410 ;
        RECT 97.060 14.990 97.520 15.180 ;
        RECT 99.920 14.990 100.370 15.180 ;
        RECT 97.060 14.760 100.370 14.990 ;
        RECT 97.060 14.680 97.520 14.760 ;
        RECT 99.920 14.670 100.370 14.760 ;
        RECT 103.760 15.410 104.210 15.500 ;
        RECT 106.610 15.410 107.070 15.490 ;
        RECT 103.760 15.180 107.070 15.410 ;
        RECT 103.760 14.990 104.210 15.180 ;
        RECT 106.610 14.990 107.070 15.180 ;
        RECT 103.760 14.760 107.070 14.990 ;
        RECT 103.760 14.670 104.210 14.760 ;
        RECT 106.610 14.680 107.070 14.760 ;
        RECT 110.560 15.410 111.020 15.490 ;
        RECT 113.420 15.410 113.870 15.500 ;
        RECT 110.560 15.180 113.870 15.410 ;
        RECT 110.560 14.990 111.020 15.180 ;
        RECT 113.420 14.990 113.870 15.180 ;
        RECT 110.560 14.760 113.870 14.990 ;
        RECT 110.560 14.680 111.020 14.760 ;
        RECT 113.420 14.670 113.870 14.760 ;
        RECT 117.260 15.410 117.710 15.500 ;
        RECT 120.110 15.410 120.570 15.490 ;
        RECT 117.260 15.180 120.570 15.410 ;
        RECT 117.260 14.990 117.710 15.180 ;
        RECT 120.110 14.990 120.570 15.180 ;
        RECT 117.260 14.760 120.570 14.990 ;
        RECT 117.260 14.670 117.710 14.760 ;
        RECT 120.110 14.680 120.570 14.760 ;
        RECT 124.060 15.410 124.520 15.490 ;
        RECT 126.920 15.410 127.370 15.500 ;
        RECT 124.060 15.180 127.370 15.410 ;
        RECT 124.060 14.990 124.520 15.180 ;
        RECT 126.920 14.990 127.370 15.180 ;
        RECT 124.060 14.760 127.370 14.990 ;
        RECT 124.060 14.680 124.520 14.760 ;
        RECT 126.920 14.670 127.370 14.760 ;
        RECT 130.760 15.410 131.210 15.500 ;
        RECT 133.610 15.410 134.070 15.490 ;
        RECT 130.760 15.180 134.070 15.410 ;
        RECT 130.760 14.990 131.210 15.180 ;
        RECT 133.610 14.990 134.070 15.180 ;
        RECT 130.760 14.760 134.070 14.990 ;
        RECT 130.760 14.670 131.210 14.760 ;
        RECT 133.610 14.680 134.070 14.760 ;
        RECT 137.560 15.410 138.020 15.490 ;
        RECT 140.420 15.410 140.870 15.500 ;
        RECT 137.560 15.180 140.870 15.410 ;
        RECT 137.560 14.990 138.020 15.180 ;
        RECT 140.420 14.990 140.870 15.180 ;
        RECT 137.560 14.760 140.870 14.990 ;
        RECT 137.560 14.680 138.020 14.760 ;
        RECT 140.420 14.670 140.870 14.760 ;
        RECT 144.260 15.410 144.710 15.500 ;
        RECT 147.110 15.410 147.570 15.490 ;
        RECT 144.260 15.180 147.570 15.410 ;
        RECT 144.260 14.990 144.710 15.180 ;
        RECT 147.110 14.990 147.570 15.180 ;
        RECT 144.260 14.760 147.570 14.990 ;
        RECT 144.260 14.670 144.710 14.760 ;
        RECT 147.110 14.680 147.570 14.760 ;
        RECT 151.060 15.410 151.520 15.490 ;
        RECT 153.920 15.410 154.370 15.500 ;
        RECT 151.060 15.180 154.370 15.410 ;
        RECT 151.060 14.990 151.520 15.180 ;
        RECT 153.920 14.990 154.370 15.180 ;
        RECT 151.060 14.760 154.370 14.990 ;
        RECT 151.060 14.680 151.520 14.760 ;
        RECT 153.920 14.670 154.370 14.760 ;
        RECT 157.760 15.410 158.210 15.500 ;
        RECT 160.610 15.410 161.070 15.490 ;
        RECT 157.760 15.180 161.070 15.410 ;
        RECT 157.760 14.990 158.210 15.180 ;
        RECT 160.610 14.990 161.070 15.180 ;
        RECT 157.760 14.760 161.070 14.990 ;
        RECT 157.760 14.670 158.210 14.760 ;
        RECT 160.610 14.680 161.070 14.760 ;
        RECT 164.560 15.410 165.020 15.490 ;
        RECT 167.420 15.410 167.870 15.500 ;
        RECT 164.560 15.180 167.870 15.410 ;
        RECT 164.560 14.990 165.020 15.180 ;
        RECT 167.420 14.990 167.870 15.180 ;
        RECT 164.560 14.760 167.870 14.990 ;
        RECT 164.560 14.680 165.020 14.760 ;
        RECT 167.420 14.670 167.870 14.760 ;
        RECT 171.260 15.410 171.710 15.500 ;
        RECT 174.110 15.410 174.570 15.490 ;
        RECT 171.260 15.180 174.570 15.410 ;
        RECT 171.260 14.990 171.710 15.180 ;
        RECT 174.110 14.990 174.570 15.180 ;
        RECT 171.260 14.760 174.570 14.990 ;
        RECT 171.260 14.670 171.710 14.760 ;
        RECT 174.110 14.680 174.570 14.760 ;
        RECT 178.060 15.410 178.520 15.490 ;
        RECT 180.920 15.410 181.370 15.500 ;
        RECT 178.060 15.180 181.370 15.410 ;
        RECT 178.060 14.990 178.520 15.180 ;
        RECT 180.920 14.990 181.370 15.180 ;
        RECT 178.060 14.760 181.370 14.990 ;
        RECT 178.060 14.680 178.520 14.760 ;
        RECT 180.920 14.670 181.370 14.760 ;
        RECT 184.760 15.410 185.210 15.500 ;
        RECT 187.610 15.410 188.070 15.490 ;
        RECT 184.760 15.180 188.070 15.410 ;
        RECT 184.760 14.990 185.210 15.180 ;
        RECT 187.610 14.990 188.070 15.180 ;
        RECT 184.760 14.760 188.070 14.990 ;
        RECT 184.760 14.670 185.210 14.760 ;
        RECT 187.610 14.680 188.070 14.760 ;
        RECT 191.560 15.410 192.020 15.490 ;
        RECT 194.420 15.410 194.870 15.500 ;
        RECT 191.560 15.180 194.870 15.410 ;
        RECT 191.560 14.990 192.020 15.180 ;
        RECT 194.420 14.990 194.870 15.180 ;
        RECT 191.560 14.760 194.870 14.990 ;
        RECT 191.560 14.680 192.020 14.760 ;
        RECT 194.420 14.670 194.870 14.760 ;
        RECT 198.260 15.410 198.710 15.500 ;
        RECT 201.110 15.410 201.570 15.490 ;
        RECT 198.260 15.180 201.570 15.410 ;
        RECT 198.260 14.990 198.710 15.180 ;
        RECT 201.110 14.990 201.570 15.180 ;
        RECT 198.260 14.760 201.570 14.990 ;
        RECT 198.260 14.670 198.710 14.760 ;
        RECT 201.110 14.680 201.570 14.760 ;
        RECT 205.060 15.410 205.520 15.490 ;
        RECT 207.920 15.410 208.370 15.500 ;
        RECT 205.060 15.180 208.370 15.410 ;
        RECT 205.060 14.990 205.520 15.180 ;
        RECT 207.920 14.990 208.370 15.180 ;
        RECT 205.060 14.760 208.370 14.990 ;
        RECT 205.060 14.680 205.520 14.760 ;
        RECT 207.920 14.670 208.370 14.760 ;
        RECT 211.760 15.410 212.210 15.500 ;
        RECT 214.610 15.410 215.070 15.490 ;
        RECT 211.760 15.180 215.070 15.410 ;
        RECT 211.760 14.990 212.210 15.180 ;
        RECT 214.610 14.990 215.070 15.180 ;
        RECT 211.760 14.760 215.070 14.990 ;
        RECT 211.760 14.670 212.210 14.760 ;
        RECT 214.610 14.680 215.070 14.760 ;
        RECT 9.260 11.800 9.710 11.890 ;
        RECT 12.110 11.800 12.570 11.880 ;
        RECT 9.260 11.570 12.570 11.800 ;
        RECT 9.260 11.380 9.710 11.570 ;
        RECT 12.110 11.380 12.570 11.570 ;
        RECT 9.260 11.150 12.570 11.380 ;
        RECT 9.260 11.060 9.710 11.150 ;
        RECT 12.110 11.070 12.570 11.150 ;
        RECT 16.060 11.800 16.520 11.880 ;
        RECT 18.920 11.800 19.370 11.890 ;
        RECT 16.060 11.570 19.370 11.800 ;
        RECT 16.060 11.380 16.520 11.570 ;
        RECT 18.920 11.380 19.370 11.570 ;
        RECT 16.060 11.150 19.370 11.380 ;
        RECT 16.060 11.070 16.520 11.150 ;
        RECT 18.920 11.060 19.370 11.150 ;
        RECT 22.760 11.800 23.210 11.890 ;
        RECT 25.610 11.800 26.070 11.880 ;
        RECT 22.760 11.570 26.070 11.800 ;
        RECT 22.760 11.380 23.210 11.570 ;
        RECT 25.610 11.380 26.070 11.570 ;
        RECT 22.760 11.150 26.070 11.380 ;
        RECT 22.760 11.060 23.210 11.150 ;
        RECT 25.610 11.070 26.070 11.150 ;
        RECT 29.560 11.800 30.020 11.880 ;
        RECT 32.420 11.800 32.870 11.890 ;
        RECT 29.560 11.570 32.870 11.800 ;
        RECT 29.560 11.380 30.020 11.570 ;
        RECT 32.420 11.380 32.870 11.570 ;
        RECT 29.560 11.150 32.870 11.380 ;
        RECT 29.560 11.070 30.020 11.150 ;
        RECT 32.420 11.060 32.870 11.150 ;
        RECT 36.260 11.800 36.710 11.890 ;
        RECT 39.110 11.800 39.570 11.880 ;
        RECT 36.260 11.570 39.570 11.800 ;
        RECT 36.260 11.380 36.710 11.570 ;
        RECT 39.110 11.380 39.570 11.570 ;
        RECT 36.260 11.150 39.570 11.380 ;
        RECT 36.260 11.060 36.710 11.150 ;
        RECT 39.110 11.070 39.570 11.150 ;
        RECT 43.060 11.800 43.520 11.880 ;
        RECT 45.920 11.800 46.370 11.890 ;
        RECT 43.060 11.570 46.370 11.800 ;
        RECT 43.060 11.380 43.520 11.570 ;
        RECT 45.920 11.380 46.370 11.570 ;
        RECT 43.060 11.150 46.370 11.380 ;
        RECT 43.060 11.070 43.520 11.150 ;
        RECT 45.920 11.060 46.370 11.150 ;
        RECT 49.760 11.800 50.210 11.890 ;
        RECT 52.610 11.800 53.070 11.880 ;
        RECT 49.760 11.570 53.070 11.800 ;
        RECT 49.760 11.380 50.210 11.570 ;
        RECT 52.610 11.380 53.070 11.570 ;
        RECT 49.760 11.150 53.070 11.380 ;
        RECT 49.760 11.060 50.210 11.150 ;
        RECT 52.610 11.070 53.070 11.150 ;
        RECT 56.560 11.800 57.020 11.880 ;
        RECT 59.420 11.800 59.870 11.890 ;
        RECT 56.560 11.570 59.870 11.800 ;
        RECT 56.560 11.380 57.020 11.570 ;
        RECT 59.420 11.380 59.870 11.570 ;
        RECT 56.560 11.150 59.870 11.380 ;
        RECT 56.560 11.070 57.020 11.150 ;
        RECT 59.420 11.060 59.870 11.150 ;
        RECT 63.260 11.800 63.710 11.890 ;
        RECT 66.110 11.800 66.570 11.880 ;
        RECT 63.260 11.570 66.570 11.800 ;
        RECT 63.260 11.380 63.710 11.570 ;
        RECT 66.110 11.380 66.570 11.570 ;
        RECT 63.260 11.150 66.570 11.380 ;
        RECT 63.260 11.060 63.710 11.150 ;
        RECT 66.110 11.070 66.570 11.150 ;
        RECT 70.060 11.800 70.520 11.880 ;
        RECT 72.920 11.800 73.370 11.890 ;
        RECT 70.060 11.570 73.370 11.800 ;
        RECT 70.060 11.380 70.520 11.570 ;
        RECT 72.920 11.380 73.370 11.570 ;
        RECT 70.060 11.150 73.370 11.380 ;
        RECT 70.060 11.070 70.520 11.150 ;
        RECT 72.920 11.060 73.370 11.150 ;
        RECT 76.760 11.800 77.210 11.890 ;
        RECT 79.610 11.800 80.070 11.880 ;
        RECT 76.760 11.570 80.070 11.800 ;
        RECT 76.760 11.380 77.210 11.570 ;
        RECT 79.610 11.380 80.070 11.570 ;
        RECT 76.760 11.150 80.070 11.380 ;
        RECT 76.760 11.060 77.210 11.150 ;
        RECT 79.610 11.070 80.070 11.150 ;
        RECT 83.560 11.800 84.020 11.880 ;
        RECT 86.420 11.800 86.870 11.890 ;
        RECT 83.560 11.570 86.870 11.800 ;
        RECT 83.560 11.380 84.020 11.570 ;
        RECT 86.420 11.380 86.870 11.570 ;
        RECT 83.560 11.150 86.870 11.380 ;
        RECT 83.560 11.070 84.020 11.150 ;
        RECT 86.420 11.060 86.870 11.150 ;
        RECT 90.260 11.800 90.710 11.890 ;
        RECT 93.110 11.800 93.570 11.880 ;
        RECT 90.260 11.570 93.570 11.800 ;
        RECT 90.260 11.380 90.710 11.570 ;
        RECT 93.110 11.380 93.570 11.570 ;
        RECT 90.260 11.150 93.570 11.380 ;
        RECT 90.260 11.060 90.710 11.150 ;
        RECT 93.110 11.070 93.570 11.150 ;
        RECT 97.060 11.800 97.520 11.880 ;
        RECT 99.920 11.800 100.370 11.890 ;
        RECT 97.060 11.570 100.370 11.800 ;
        RECT 97.060 11.380 97.520 11.570 ;
        RECT 99.920 11.380 100.370 11.570 ;
        RECT 97.060 11.150 100.370 11.380 ;
        RECT 97.060 11.070 97.520 11.150 ;
        RECT 99.920 11.060 100.370 11.150 ;
        RECT 103.760 11.800 104.210 11.890 ;
        RECT 106.610 11.800 107.070 11.880 ;
        RECT 103.760 11.570 107.070 11.800 ;
        RECT 103.760 11.380 104.210 11.570 ;
        RECT 106.610 11.380 107.070 11.570 ;
        RECT 103.760 11.150 107.070 11.380 ;
        RECT 103.760 11.060 104.210 11.150 ;
        RECT 106.610 11.070 107.070 11.150 ;
        RECT 110.560 11.800 111.020 11.880 ;
        RECT 113.420 11.800 113.870 11.890 ;
        RECT 110.560 11.570 113.870 11.800 ;
        RECT 110.560 11.380 111.020 11.570 ;
        RECT 113.420 11.380 113.870 11.570 ;
        RECT 110.560 11.150 113.870 11.380 ;
        RECT 110.560 11.070 111.020 11.150 ;
        RECT 113.420 11.060 113.870 11.150 ;
        RECT 117.260 11.800 117.710 11.890 ;
        RECT 120.110 11.800 120.570 11.880 ;
        RECT 117.260 11.570 120.570 11.800 ;
        RECT 117.260 11.380 117.710 11.570 ;
        RECT 120.110 11.380 120.570 11.570 ;
        RECT 117.260 11.150 120.570 11.380 ;
        RECT 117.260 11.060 117.710 11.150 ;
        RECT 120.110 11.070 120.570 11.150 ;
        RECT 124.060 11.800 124.520 11.880 ;
        RECT 126.920 11.800 127.370 11.890 ;
        RECT 124.060 11.570 127.370 11.800 ;
        RECT 124.060 11.380 124.520 11.570 ;
        RECT 126.920 11.380 127.370 11.570 ;
        RECT 124.060 11.150 127.370 11.380 ;
        RECT 124.060 11.070 124.520 11.150 ;
        RECT 126.920 11.060 127.370 11.150 ;
        RECT 130.760 11.800 131.210 11.890 ;
        RECT 133.610 11.800 134.070 11.880 ;
        RECT 130.760 11.570 134.070 11.800 ;
        RECT 130.760 11.380 131.210 11.570 ;
        RECT 133.610 11.380 134.070 11.570 ;
        RECT 130.760 11.150 134.070 11.380 ;
        RECT 130.760 11.060 131.210 11.150 ;
        RECT 133.610 11.070 134.070 11.150 ;
        RECT 137.560 11.800 138.020 11.880 ;
        RECT 140.420 11.800 140.870 11.890 ;
        RECT 137.560 11.570 140.870 11.800 ;
        RECT 137.560 11.380 138.020 11.570 ;
        RECT 140.420 11.380 140.870 11.570 ;
        RECT 137.560 11.150 140.870 11.380 ;
        RECT 137.560 11.070 138.020 11.150 ;
        RECT 140.420 11.060 140.870 11.150 ;
        RECT 144.260 11.800 144.710 11.890 ;
        RECT 147.110 11.800 147.570 11.880 ;
        RECT 144.260 11.570 147.570 11.800 ;
        RECT 144.260 11.380 144.710 11.570 ;
        RECT 147.110 11.380 147.570 11.570 ;
        RECT 144.260 11.150 147.570 11.380 ;
        RECT 144.260 11.060 144.710 11.150 ;
        RECT 147.110 11.070 147.570 11.150 ;
        RECT 151.060 11.800 151.520 11.880 ;
        RECT 153.920 11.800 154.370 11.890 ;
        RECT 151.060 11.570 154.370 11.800 ;
        RECT 151.060 11.380 151.520 11.570 ;
        RECT 153.920 11.380 154.370 11.570 ;
        RECT 151.060 11.150 154.370 11.380 ;
        RECT 151.060 11.070 151.520 11.150 ;
        RECT 153.920 11.060 154.370 11.150 ;
        RECT 157.760 11.800 158.210 11.890 ;
        RECT 160.610 11.800 161.070 11.880 ;
        RECT 157.760 11.570 161.070 11.800 ;
        RECT 157.760 11.380 158.210 11.570 ;
        RECT 160.610 11.380 161.070 11.570 ;
        RECT 157.760 11.150 161.070 11.380 ;
        RECT 157.760 11.060 158.210 11.150 ;
        RECT 160.610 11.070 161.070 11.150 ;
        RECT 164.560 11.800 165.020 11.880 ;
        RECT 167.420 11.800 167.870 11.890 ;
        RECT 164.560 11.570 167.870 11.800 ;
        RECT 164.560 11.380 165.020 11.570 ;
        RECT 167.420 11.380 167.870 11.570 ;
        RECT 164.560 11.150 167.870 11.380 ;
        RECT 164.560 11.070 165.020 11.150 ;
        RECT 167.420 11.060 167.870 11.150 ;
        RECT 171.260 11.800 171.710 11.890 ;
        RECT 174.110 11.800 174.570 11.880 ;
        RECT 171.260 11.570 174.570 11.800 ;
        RECT 171.260 11.380 171.710 11.570 ;
        RECT 174.110 11.380 174.570 11.570 ;
        RECT 171.260 11.150 174.570 11.380 ;
        RECT 171.260 11.060 171.710 11.150 ;
        RECT 174.110 11.070 174.570 11.150 ;
        RECT 178.060 11.800 178.520 11.880 ;
        RECT 180.920 11.800 181.370 11.890 ;
        RECT 178.060 11.570 181.370 11.800 ;
        RECT 178.060 11.380 178.520 11.570 ;
        RECT 180.920 11.380 181.370 11.570 ;
        RECT 178.060 11.150 181.370 11.380 ;
        RECT 178.060 11.070 178.520 11.150 ;
        RECT 180.920 11.060 181.370 11.150 ;
        RECT 184.760 11.800 185.210 11.890 ;
        RECT 187.610 11.800 188.070 11.880 ;
        RECT 184.760 11.570 188.070 11.800 ;
        RECT 184.760 11.380 185.210 11.570 ;
        RECT 187.610 11.380 188.070 11.570 ;
        RECT 184.760 11.150 188.070 11.380 ;
        RECT 184.760 11.060 185.210 11.150 ;
        RECT 187.610 11.070 188.070 11.150 ;
        RECT 191.560 11.800 192.020 11.880 ;
        RECT 194.420 11.800 194.870 11.890 ;
        RECT 191.560 11.570 194.870 11.800 ;
        RECT 191.560 11.380 192.020 11.570 ;
        RECT 194.420 11.380 194.870 11.570 ;
        RECT 191.560 11.150 194.870 11.380 ;
        RECT 191.560 11.070 192.020 11.150 ;
        RECT 194.420 11.060 194.870 11.150 ;
        RECT 198.260 11.800 198.710 11.890 ;
        RECT 201.110 11.800 201.570 11.880 ;
        RECT 198.260 11.570 201.570 11.800 ;
        RECT 198.260 11.380 198.710 11.570 ;
        RECT 201.110 11.380 201.570 11.570 ;
        RECT 198.260 11.150 201.570 11.380 ;
        RECT 198.260 11.060 198.710 11.150 ;
        RECT 201.110 11.070 201.570 11.150 ;
        RECT 205.060 11.800 205.520 11.880 ;
        RECT 207.920 11.800 208.370 11.890 ;
        RECT 205.060 11.570 208.370 11.800 ;
        RECT 205.060 11.380 205.520 11.570 ;
        RECT 207.920 11.380 208.370 11.570 ;
        RECT 205.060 11.150 208.370 11.380 ;
        RECT 205.060 11.070 205.520 11.150 ;
        RECT 207.920 11.060 208.370 11.150 ;
        RECT 211.760 11.800 212.210 11.890 ;
        RECT 214.610 11.800 215.070 11.880 ;
        RECT 211.760 11.570 215.070 11.800 ;
        RECT 211.760 11.380 212.210 11.570 ;
        RECT 214.610 11.380 215.070 11.570 ;
        RECT 211.760 11.150 215.070 11.380 ;
        RECT 211.760 11.060 212.210 11.150 ;
        RECT 214.610 11.070 215.070 11.150 ;
        RECT 9.260 8.190 9.710 8.280 ;
        RECT 12.110 8.190 12.570 8.270 ;
        RECT 9.260 7.960 12.570 8.190 ;
        RECT 9.260 7.770 9.710 7.960 ;
        RECT 12.110 7.770 12.570 7.960 ;
        RECT 9.260 7.540 12.570 7.770 ;
        RECT 9.260 7.450 9.710 7.540 ;
        RECT 12.110 7.460 12.570 7.540 ;
        RECT 16.060 8.190 16.520 8.270 ;
        RECT 18.920 8.190 19.370 8.280 ;
        RECT 16.060 7.960 19.370 8.190 ;
        RECT 16.060 7.770 16.520 7.960 ;
        RECT 18.920 7.770 19.370 7.960 ;
        RECT 16.060 7.540 19.370 7.770 ;
        RECT 16.060 7.460 16.520 7.540 ;
        RECT 18.920 7.450 19.370 7.540 ;
        RECT 22.760 8.190 23.210 8.280 ;
        RECT 25.610 8.190 26.070 8.270 ;
        RECT 22.760 7.960 26.070 8.190 ;
        RECT 22.760 7.770 23.210 7.960 ;
        RECT 25.610 7.770 26.070 7.960 ;
        RECT 22.760 7.540 26.070 7.770 ;
        RECT 22.760 7.450 23.210 7.540 ;
        RECT 25.610 7.460 26.070 7.540 ;
        RECT 29.560 8.190 30.020 8.270 ;
        RECT 32.420 8.190 32.870 8.280 ;
        RECT 29.560 7.960 32.870 8.190 ;
        RECT 29.560 7.770 30.020 7.960 ;
        RECT 32.420 7.770 32.870 7.960 ;
        RECT 29.560 7.540 32.870 7.770 ;
        RECT 29.560 7.460 30.020 7.540 ;
        RECT 32.420 7.450 32.870 7.540 ;
        RECT 36.260 8.190 36.710 8.280 ;
        RECT 39.110 8.190 39.570 8.270 ;
        RECT 36.260 7.960 39.570 8.190 ;
        RECT 36.260 7.770 36.710 7.960 ;
        RECT 39.110 7.770 39.570 7.960 ;
        RECT 36.260 7.540 39.570 7.770 ;
        RECT 36.260 7.450 36.710 7.540 ;
        RECT 39.110 7.460 39.570 7.540 ;
        RECT 43.060 8.190 43.520 8.270 ;
        RECT 45.920 8.190 46.370 8.280 ;
        RECT 43.060 7.960 46.370 8.190 ;
        RECT 43.060 7.770 43.520 7.960 ;
        RECT 45.920 7.770 46.370 7.960 ;
        RECT 43.060 7.540 46.370 7.770 ;
        RECT 43.060 7.460 43.520 7.540 ;
        RECT 45.920 7.450 46.370 7.540 ;
        RECT 49.760 8.190 50.210 8.280 ;
        RECT 52.610 8.190 53.070 8.270 ;
        RECT 49.760 7.960 53.070 8.190 ;
        RECT 49.760 7.770 50.210 7.960 ;
        RECT 52.610 7.770 53.070 7.960 ;
        RECT 49.760 7.540 53.070 7.770 ;
        RECT 49.760 7.450 50.210 7.540 ;
        RECT 52.610 7.460 53.070 7.540 ;
        RECT 56.560 8.190 57.020 8.270 ;
        RECT 59.420 8.190 59.870 8.280 ;
        RECT 56.560 7.960 59.870 8.190 ;
        RECT 56.560 7.770 57.020 7.960 ;
        RECT 59.420 7.770 59.870 7.960 ;
        RECT 56.560 7.540 59.870 7.770 ;
        RECT 56.560 7.460 57.020 7.540 ;
        RECT 59.420 7.450 59.870 7.540 ;
        RECT 63.260 8.190 63.710 8.280 ;
        RECT 66.110 8.190 66.570 8.270 ;
        RECT 63.260 7.960 66.570 8.190 ;
        RECT 63.260 7.770 63.710 7.960 ;
        RECT 66.110 7.770 66.570 7.960 ;
        RECT 63.260 7.540 66.570 7.770 ;
        RECT 63.260 7.450 63.710 7.540 ;
        RECT 66.110 7.460 66.570 7.540 ;
        RECT 70.060 8.190 70.520 8.270 ;
        RECT 72.920 8.190 73.370 8.280 ;
        RECT 70.060 7.960 73.370 8.190 ;
        RECT 70.060 7.770 70.520 7.960 ;
        RECT 72.920 7.770 73.370 7.960 ;
        RECT 70.060 7.540 73.370 7.770 ;
        RECT 70.060 7.460 70.520 7.540 ;
        RECT 72.920 7.450 73.370 7.540 ;
        RECT 76.760 8.190 77.210 8.280 ;
        RECT 79.610 8.190 80.070 8.270 ;
        RECT 76.760 7.960 80.070 8.190 ;
        RECT 76.760 7.770 77.210 7.960 ;
        RECT 79.610 7.770 80.070 7.960 ;
        RECT 76.760 7.540 80.070 7.770 ;
        RECT 76.760 7.450 77.210 7.540 ;
        RECT 79.610 7.460 80.070 7.540 ;
        RECT 83.560 8.190 84.020 8.270 ;
        RECT 86.420 8.190 86.870 8.280 ;
        RECT 83.560 7.960 86.870 8.190 ;
        RECT 83.560 7.770 84.020 7.960 ;
        RECT 86.420 7.770 86.870 7.960 ;
        RECT 83.560 7.540 86.870 7.770 ;
        RECT 83.560 7.460 84.020 7.540 ;
        RECT 86.420 7.450 86.870 7.540 ;
        RECT 90.260 8.190 90.710 8.280 ;
        RECT 93.110 8.190 93.570 8.270 ;
        RECT 90.260 7.960 93.570 8.190 ;
        RECT 90.260 7.770 90.710 7.960 ;
        RECT 93.110 7.770 93.570 7.960 ;
        RECT 90.260 7.540 93.570 7.770 ;
        RECT 90.260 7.450 90.710 7.540 ;
        RECT 93.110 7.460 93.570 7.540 ;
        RECT 97.060 8.190 97.520 8.270 ;
        RECT 99.920 8.190 100.370 8.280 ;
        RECT 97.060 7.960 100.370 8.190 ;
        RECT 97.060 7.770 97.520 7.960 ;
        RECT 99.920 7.770 100.370 7.960 ;
        RECT 97.060 7.540 100.370 7.770 ;
        RECT 97.060 7.460 97.520 7.540 ;
        RECT 99.920 7.450 100.370 7.540 ;
        RECT 103.760 8.190 104.210 8.280 ;
        RECT 106.610 8.190 107.070 8.270 ;
        RECT 103.760 7.960 107.070 8.190 ;
        RECT 103.760 7.770 104.210 7.960 ;
        RECT 106.610 7.770 107.070 7.960 ;
        RECT 103.760 7.540 107.070 7.770 ;
        RECT 103.760 7.450 104.210 7.540 ;
        RECT 106.610 7.460 107.070 7.540 ;
        RECT 110.560 8.190 111.020 8.270 ;
        RECT 113.420 8.190 113.870 8.280 ;
        RECT 110.560 7.960 113.870 8.190 ;
        RECT 110.560 7.770 111.020 7.960 ;
        RECT 113.420 7.770 113.870 7.960 ;
        RECT 110.560 7.540 113.870 7.770 ;
        RECT 110.560 7.460 111.020 7.540 ;
        RECT 113.420 7.450 113.870 7.540 ;
        RECT 117.260 8.190 117.710 8.280 ;
        RECT 120.110 8.190 120.570 8.270 ;
        RECT 117.260 7.960 120.570 8.190 ;
        RECT 117.260 7.770 117.710 7.960 ;
        RECT 120.110 7.770 120.570 7.960 ;
        RECT 117.260 7.540 120.570 7.770 ;
        RECT 117.260 7.450 117.710 7.540 ;
        RECT 120.110 7.460 120.570 7.540 ;
        RECT 124.060 8.190 124.520 8.270 ;
        RECT 126.920 8.190 127.370 8.280 ;
        RECT 124.060 7.960 127.370 8.190 ;
        RECT 124.060 7.770 124.520 7.960 ;
        RECT 126.920 7.770 127.370 7.960 ;
        RECT 124.060 7.540 127.370 7.770 ;
        RECT 124.060 7.460 124.520 7.540 ;
        RECT 126.920 7.450 127.370 7.540 ;
        RECT 130.760 8.190 131.210 8.280 ;
        RECT 133.610 8.190 134.070 8.270 ;
        RECT 130.760 7.960 134.070 8.190 ;
        RECT 130.760 7.770 131.210 7.960 ;
        RECT 133.610 7.770 134.070 7.960 ;
        RECT 130.760 7.540 134.070 7.770 ;
        RECT 130.760 7.450 131.210 7.540 ;
        RECT 133.610 7.460 134.070 7.540 ;
        RECT 137.560 8.190 138.020 8.270 ;
        RECT 140.420 8.190 140.870 8.280 ;
        RECT 137.560 7.960 140.870 8.190 ;
        RECT 137.560 7.770 138.020 7.960 ;
        RECT 140.420 7.770 140.870 7.960 ;
        RECT 137.560 7.540 140.870 7.770 ;
        RECT 137.560 7.460 138.020 7.540 ;
        RECT 140.420 7.450 140.870 7.540 ;
        RECT 144.260 8.190 144.710 8.280 ;
        RECT 147.110 8.190 147.570 8.270 ;
        RECT 144.260 7.960 147.570 8.190 ;
        RECT 144.260 7.770 144.710 7.960 ;
        RECT 147.110 7.770 147.570 7.960 ;
        RECT 144.260 7.540 147.570 7.770 ;
        RECT 144.260 7.450 144.710 7.540 ;
        RECT 147.110 7.460 147.570 7.540 ;
        RECT 151.060 8.190 151.520 8.270 ;
        RECT 153.920 8.190 154.370 8.280 ;
        RECT 151.060 7.960 154.370 8.190 ;
        RECT 151.060 7.770 151.520 7.960 ;
        RECT 153.920 7.770 154.370 7.960 ;
        RECT 151.060 7.540 154.370 7.770 ;
        RECT 151.060 7.460 151.520 7.540 ;
        RECT 153.920 7.450 154.370 7.540 ;
        RECT 157.760 8.190 158.210 8.280 ;
        RECT 160.610 8.190 161.070 8.270 ;
        RECT 157.760 7.960 161.070 8.190 ;
        RECT 157.760 7.770 158.210 7.960 ;
        RECT 160.610 7.770 161.070 7.960 ;
        RECT 157.760 7.540 161.070 7.770 ;
        RECT 157.760 7.450 158.210 7.540 ;
        RECT 160.610 7.460 161.070 7.540 ;
        RECT 164.560 8.190 165.020 8.270 ;
        RECT 167.420 8.190 167.870 8.280 ;
        RECT 164.560 7.960 167.870 8.190 ;
        RECT 164.560 7.770 165.020 7.960 ;
        RECT 167.420 7.770 167.870 7.960 ;
        RECT 164.560 7.540 167.870 7.770 ;
        RECT 164.560 7.460 165.020 7.540 ;
        RECT 167.420 7.450 167.870 7.540 ;
        RECT 171.260 8.190 171.710 8.280 ;
        RECT 174.110 8.190 174.570 8.270 ;
        RECT 171.260 7.960 174.570 8.190 ;
        RECT 171.260 7.770 171.710 7.960 ;
        RECT 174.110 7.770 174.570 7.960 ;
        RECT 171.260 7.540 174.570 7.770 ;
        RECT 171.260 7.450 171.710 7.540 ;
        RECT 174.110 7.460 174.570 7.540 ;
        RECT 178.060 8.190 178.520 8.270 ;
        RECT 180.920 8.190 181.370 8.280 ;
        RECT 178.060 7.960 181.370 8.190 ;
        RECT 178.060 7.770 178.520 7.960 ;
        RECT 180.920 7.770 181.370 7.960 ;
        RECT 178.060 7.540 181.370 7.770 ;
        RECT 178.060 7.460 178.520 7.540 ;
        RECT 180.920 7.450 181.370 7.540 ;
        RECT 184.760 8.190 185.210 8.280 ;
        RECT 187.610 8.190 188.070 8.270 ;
        RECT 184.760 7.960 188.070 8.190 ;
        RECT 184.760 7.770 185.210 7.960 ;
        RECT 187.610 7.770 188.070 7.960 ;
        RECT 184.760 7.540 188.070 7.770 ;
        RECT 184.760 7.450 185.210 7.540 ;
        RECT 187.610 7.460 188.070 7.540 ;
        RECT 191.560 8.190 192.020 8.270 ;
        RECT 194.420 8.190 194.870 8.280 ;
        RECT 191.560 7.960 194.870 8.190 ;
        RECT 191.560 7.770 192.020 7.960 ;
        RECT 194.420 7.770 194.870 7.960 ;
        RECT 191.560 7.540 194.870 7.770 ;
        RECT 191.560 7.460 192.020 7.540 ;
        RECT 194.420 7.450 194.870 7.540 ;
        RECT 198.260 8.190 198.710 8.280 ;
        RECT 201.110 8.190 201.570 8.270 ;
        RECT 198.260 7.960 201.570 8.190 ;
        RECT 198.260 7.770 198.710 7.960 ;
        RECT 201.110 7.770 201.570 7.960 ;
        RECT 198.260 7.540 201.570 7.770 ;
        RECT 198.260 7.450 198.710 7.540 ;
        RECT 201.110 7.460 201.570 7.540 ;
        RECT 205.060 8.190 205.520 8.270 ;
        RECT 207.920 8.190 208.370 8.280 ;
        RECT 205.060 7.960 208.370 8.190 ;
        RECT 205.060 7.770 205.520 7.960 ;
        RECT 207.920 7.770 208.370 7.960 ;
        RECT 205.060 7.540 208.370 7.770 ;
        RECT 205.060 7.460 205.520 7.540 ;
        RECT 207.920 7.450 208.370 7.540 ;
        RECT 211.760 8.190 212.210 8.280 ;
        RECT 214.610 8.190 215.070 8.270 ;
        RECT 211.760 7.960 215.070 8.190 ;
        RECT 211.760 7.770 212.210 7.960 ;
        RECT 214.610 7.770 215.070 7.960 ;
        RECT 211.760 7.540 215.070 7.770 ;
        RECT 211.760 7.450 212.210 7.540 ;
        RECT 214.610 7.460 215.070 7.540 ;
        RECT 9.260 4.580 9.710 4.670 ;
        RECT 12.110 4.580 12.570 4.660 ;
        RECT 9.260 4.350 12.570 4.580 ;
        RECT 9.260 4.160 9.710 4.350 ;
        RECT 12.110 4.160 12.570 4.350 ;
        RECT 9.260 3.930 12.570 4.160 ;
        RECT 9.260 3.840 9.710 3.930 ;
        RECT 12.110 3.850 12.570 3.930 ;
        RECT 16.060 4.580 16.520 4.660 ;
        RECT 18.920 4.580 19.370 4.670 ;
        RECT 16.060 4.350 19.370 4.580 ;
        RECT 16.060 4.160 16.520 4.350 ;
        RECT 18.920 4.160 19.370 4.350 ;
        RECT 16.060 3.930 19.370 4.160 ;
        RECT 16.060 3.850 16.520 3.930 ;
        RECT 18.920 3.840 19.370 3.930 ;
        RECT 22.760 4.580 23.210 4.670 ;
        RECT 25.610 4.580 26.070 4.660 ;
        RECT 22.760 4.350 26.070 4.580 ;
        RECT 22.760 4.160 23.210 4.350 ;
        RECT 25.610 4.160 26.070 4.350 ;
        RECT 22.760 3.930 26.070 4.160 ;
        RECT 22.760 3.840 23.210 3.930 ;
        RECT 25.610 3.850 26.070 3.930 ;
        RECT 29.560 4.580 30.020 4.660 ;
        RECT 32.420 4.580 32.870 4.670 ;
        RECT 29.560 4.350 32.870 4.580 ;
        RECT 29.560 4.160 30.020 4.350 ;
        RECT 32.420 4.160 32.870 4.350 ;
        RECT 29.560 3.930 32.870 4.160 ;
        RECT 29.560 3.850 30.020 3.930 ;
        RECT 32.420 3.840 32.870 3.930 ;
        RECT 36.260 4.580 36.710 4.670 ;
        RECT 39.110 4.580 39.570 4.660 ;
        RECT 36.260 4.350 39.570 4.580 ;
        RECT 36.260 4.160 36.710 4.350 ;
        RECT 39.110 4.160 39.570 4.350 ;
        RECT 36.260 3.930 39.570 4.160 ;
        RECT 36.260 3.840 36.710 3.930 ;
        RECT 39.110 3.850 39.570 3.930 ;
        RECT 43.060 4.580 43.520 4.660 ;
        RECT 45.920 4.580 46.370 4.670 ;
        RECT 43.060 4.350 46.370 4.580 ;
        RECT 43.060 4.160 43.520 4.350 ;
        RECT 45.920 4.160 46.370 4.350 ;
        RECT 43.060 3.930 46.370 4.160 ;
        RECT 43.060 3.850 43.520 3.930 ;
        RECT 45.920 3.840 46.370 3.930 ;
        RECT 49.760 4.580 50.210 4.670 ;
        RECT 52.610 4.580 53.070 4.660 ;
        RECT 49.760 4.350 53.070 4.580 ;
        RECT 49.760 4.160 50.210 4.350 ;
        RECT 52.610 4.160 53.070 4.350 ;
        RECT 49.760 3.930 53.070 4.160 ;
        RECT 49.760 3.840 50.210 3.930 ;
        RECT 52.610 3.850 53.070 3.930 ;
        RECT 56.560 4.580 57.020 4.660 ;
        RECT 59.420 4.580 59.870 4.670 ;
        RECT 56.560 4.350 59.870 4.580 ;
        RECT 56.560 4.160 57.020 4.350 ;
        RECT 59.420 4.160 59.870 4.350 ;
        RECT 56.560 3.930 59.870 4.160 ;
        RECT 56.560 3.850 57.020 3.930 ;
        RECT 59.420 3.840 59.870 3.930 ;
        RECT 63.260 4.580 63.710 4.670 ;
        RECT 66.110 4.580 66.570 4.660 ;
        RECT 63.260 4.350 66.570 4.580 ;
        RECT 63.260 4.160 63.710 4.350 ;
        RECT 66.110 4.160 66.570 4.350 ;
        RECT 63.260 3.930 66.570 4.160 ;
        RECT 63.260 3.840 63.710 3.930 ;
        RECT 66.110 3.850 66.570 3.930 ;
        RECT 70.060 4.580 70.520 4.660 ;
        RECT 72.920 4.580 73.370 4.670 ;
        RECT 70.060 4.350 73.370 4.580 ;
        RECT 70.060 4.160 70.520 4.350 ;
        RECT 72.920 4.160 73.370 4.350 ;
        RECT 70.060 3.930 73.370 4.160 ;
        RECT 70.060 3.850 70.520 3.930 ;
        RECT 72.920 3.840 73.370 3.930 ;
        RECT 76.760 4.580 77.210 4.670 ;
        RECT 79.610 4.580 80.070 4.660 ;
        RECT 76.760 4.350 80.070 4.580 ;
        RECT 76.760 4.160 77.210 4.350 ;
        RECT 79.610 4.160 80.070 4.350 ;
        RECT 76.760 3.930 80.070 4.160 ;
        RECT 76.760 3.840 77.210 3.930 ;
        RECT 79.610 3.850 80.070 3.930 ;
        RECT 83.560 4.580 84.020 4.660 ;
        RECT 86.420 4.580 86.870 4.670 ;
        RECT 83.560 4.350 86.870 4.580 ;
        RECT 83.560 4.160 84.020 4.350 ;
        RECT 86.420 4.160 86.870 4.350 ;
        RECT 83.560 3.930 86.870 4.160 ;
        RECT 83.560 3.850 84.020 3.930 ;
        RECT 86.420 3.840 86.870 3.930 ;
        RECT 90.260 4.580 90.710 4.670 ;
        RECT 93.110 4.580 93.570 4.660 ;
        RECT 90.260 4.350 93.570 4.580 ;
        RECT 90.260 4.160 90.710 4.350 ;
        RECT 93.110 4.160 93.570 4.350 ;
        RECT 90.260 3.930 93.570 4.160 ;
        RECT 90.260 3.840 90.710 3.930 ;
        RECT 93.110 3.850 93.570 3.930 ;
        RECT 97.060 4.580 97.520 4.660 ;
        RECT 99.920 4.580 100.370 4.670 ;
        RECT 97.060 4.350 100.370 4.580 ;
        RECT 97.060 4.160 97.520 4.350 ;
        RECT 99.920 4.160 100.370 4.350 ;
        RECT 97.060 3.930 100.370 4.160 ;
        RECT 97.060 3.850 97.520 3.930 ;
        RECT 99.920 3.840 100.370 3.930 ;
        RECT 103.760 4.580 104.210 4.670 ;
        RECT 106.610 4.580 107.070 4.660 ;
        RECT 103.760 4.350 107.070 4.580 ;
        RECT 103.760 4.160 104.210 4.350 ;
        RECT 106.610 4.160 107.070 4.350 ;
        RECT 103.760 3.930 107.070 4.160 ;
        RECT 103.760 3.840 104.210 3.930 ;
        RECT 106.610 3.850 107.070 3.930 ;
        RECT 110.560 4.580 111.020 4.660 ;
        RECT 113.420 4.580 113.870 4.670 ;
        RECT 110.560 4.350 113.870 4.580 ;
        RECT 110.560 4.160 111.020 4.350 ;
        RECT 113.420 4.160 113.870 4.350 ;
        RECT 110.560 3.930 113.870 4.160 ;
        RECT 110.560 3.850 111.020 3.930 ;
        RECT 113.420 3.840 113.870 3.930 ;
        RECT 117.260 4.580 117.710 4.670 ;
        RECT 120.110 4.580 120.570 4.660 ;
        RECT 117.260 4.350 120.570 4.580 ;
        RECT 117.260 4.160 117.710 4.350 ;
        RECT 120.110 4.160 120.570 4.350 ;
        RECT 117.260 3.930 120.570 4.160 ;
        RECT 117.260 3.840 117.710 3.930 ;
        RECT 120.110 3.850 120.570 3.930 ;
        RECT 124.060 4.580 124.520 4.660 ;
        RECT 126.920 4.580 127.370 4.670 ;
        RECT 124.060 4.350 127.370 4.580 ;
        RECT 124.060 4.160 124.520 4.350 ;
        RECT 126.920 4.160 127.370 4.350 ;
        RECT 124.060 3.930 127.370 4.160 ;
        RECT 124.060 3.850 124.520 3.930 ;
        RECT 126.920 3.840 127.370 3.930 ;
        RECT 130.760 4.580 131.210 4.670 ;
        RECT 133.610 4.580 134.070 4.660 ;
        RECT 130.760 4.350 134.070 4.580 ;
        RECT 130.760 4.160 131.210 4.350 ;
        RECT 133.610 4.160 134.070 4.350 ;
        RECT 130.760 3.930 134.070 4.160 ;
        RECT 130.760 3.840 131.210 3.930 ;
        RECT 133.610 3.850 134.070 3.930 ;
        RECT 137.560 4.580 138.020 4.660 ;
        RECT 140.420 4.580 140.870 4.670 ;
        RECT 137.560 4.350 140.870 4.580 ;
        RECT 137.560 4.160 138.020 4.350 ;
        RECT 140.420 4.160 140.870 4.350 ;
        RECT 137.560 3.930 140.870 4.160 ;
        RECT 137.560 3.850 138.020 3.930 ;
        RECT 140.420 3.840 140.870 3.930 ;
        RECT 144.260 4.580 144.710 4.670 ;
        RECT 147.110 4.580 147.570 4.660 ;
        RECT 144.260 4.350 147.570 4.580 ;
        RECT 144.260 4.160 144.710 4.350 ;
        RECT 147.110 4.160 147.570 4.350 ;
        RECT 144.260 3.930 147.570 4.160 ;
        RECT 144.260 3.840 144.710 3.930 ;
        RECT 147.110 3.850 147.570 3.930 ;
        RECT 151.060 4.580 151.520 4.660 ;
        RECT 153.920 4.580 154.370 4.670 ;
        RECT 151.060 4.350 154.370 4.580 ;
        RECT 151.060 4.160 151.520 4.350 ;
        RECT 153.920 4.160 154.370 4.350 ;
        RECT 151.060 3.930 154.370 4.160 ;
        RECT 151.060 3.850 151.520 3.930 ;
        RECT 153.920 3.840 154.370 3.930 ;
        RECT 157.760 4.580 158.210 4.670 ;
        RECT 160.610 4.580 161.070 4.660 ;
        RECT 157.760 4.350 161.070 4.580 ;
        RECT 157.760 4.160 158.210 4.350 ;
        RECT 160.610 4.160 161.070 4.350 ;
        RECT 157.760 3.930 161.070 4.160 ;
        RECT 157.760 3.840 158.210 3.930 ;
        RECT 160.610 3.850 161.070 3.930 ;
        RECT 164.560 4.580 165.020 4.660 ;
        RECT 167.420 4.580 167.870 4.670 ;
        RECT 164.560 4.350 167.870 4.580 ;
        RECT 164.560 4.160 165.020 4.350 ;
        RECT 167.420 4.160 167.870 4.350 ;
        RECT 164.560 3.930 167.870 4.160 ;
        RECT 164.560 3.850 165.020 3.930 ;
        RECT 167.420 3.840 167.870 3.930 ;
        RECT 171.260 4.580 171.710 4.670 ;
        RECT 174.110 4.580 174.570 4.660 ;
        RECT 171.260 4.350 174.570 4.580 ;
        RECT 171.260 4.160 171.710 4.350 ;
        RECT 174.110 4.160 174.570 4.350 ;
        RECT 171.260 3.930 174.570 4.160 ;
        RECT 171.260 3.840 171.710 3.930 ;
        RECT 174.110 3.850 174.570 3.930 ;
        RECT 178.060 4.580 178.520 4.660 ;
        RECT 180.920 4.580 181.370 4.670 ;
        RECT 178.060 4.350 181.370 4.580 ;
        RECT 178.060 4.160 178.520 4.350 ;
        RECT 180.920 4.160 181.370 4.350 ;
        RECT 178.060 3.930 181.370 4.160 ;
        RECT 178.060 3.850 178.520 3.930 ;
        RECT 180.920 3.840 181.370 3.930 ;
        RECT 184.760 4.580 185.210 4.670 ;
        RECT 187.610 4.580 188.070 4.660 ;
        RECT 184.760 4.350 188.070 4.580 ;
        RECT 184.760 4.160 185.210 4.350 ;
        RECT 187.610 4.160 188.070 4.350 ;
        RECT 184.760 3.930 188.070 4.160 ;
        RECT 184.760 3.840 185.210 3.930 ;
        RECT 187.610 3.850 188.070 3.930 ;
        RECT 191.560 4.580 192.020 4.660 ;
        RECT 194.420 4.580 194.870 4.670 ;
        RECT 191.560 4.350 194.870 4.580 ;
        RECT 191.560 4.160 192.020 4.350 ;
        RECT 194.420 4.160 194.870 4.350 ;
        RECT 191.560 3.930 194.870 4.160 ;
        RECT 191.560 3.850 192.020 3.930 ;
        RECT 194.420 3.840 194.870 3.930 ;
        RECT 198.260 4.580 198.710 4.670 ;
        RECT 201.110 4.580 201.570 4.660 ;
        RECT 198.260 4.350 201.570 4.580 ;
        RECT 198.260 4.160 198.710 4.350 ;
        RECT 201.110 4.160 201.570 4.350 ;
        RECT 198.260 3.930 201.570 4.160 ;
        RECT 198.260 3.840 198.710 3.930 ;
        RECT 201.110 3.850 201.570 3.930 ;
        RECT 205.060 4.580 205.520 4.660 ;
        RECT 207.920 4.580 208.370 4.670 ;
        RECT 205.060 4.350 208.370 4.580 ;
        RECT 205.060 4.160 205.520 4.350 ;
        RECT 207.920 4.160 208.370 4.350 ;
        RECT 205.060 3.930 208.370 4.160 ;
        RECT 205.060 3.850 205.520 3.930 ;
        RECT 207.920 3.840 208.370 3.930 ;
        RECT 211.760 4.580 212.210 4.670 ;
        RECT 214.610 4.580 215.070 4.660 ;
        RECT 211.760 4.350 215.070 4.580 ;
        RECT 211.760 4.160 212.210 4.350 ;
        RECT 214.610 4.160 215.070 4.350 ;
        RECT 211.760 3.930 215.070 4.160 ;
        RECT 211.760 3.840 212.210 3.930 ;
        RECT 214.610 3.850 215.070 3.930 ;
        RECT 9.260 0.970 9.710 1.060 ;
        RECT 12.110 0.970 12.570 1.050 ;
        RECT 9.260 0.740 12.570 0.970 ;
        RECT 9.260 0.550 9.710 0.740 ;
        RECT 12.110 0.550 12.570 0.740 ;
        RECT 9.260 0.320 12.570 0.550 ;
        RECT 9.260 0.230 9.710 0.320 ;
        RECT 12.110 0.240 12.570 0.320 ;
        RECT 16.060 0.970 16.520 1.050 ;
        RECT 18.920 0.970 19.370 1.060 ;
        RECT 16.060 0.740 19.370 0.970 ;
        RECT 16.060 0.550 16.520 0.740 ;
        RECT 18.920 0.550 19.370 0.740 ;
        RECT 16.060 0.320 19.370 0.550 ;
        RECT 16.060 0.240 16.520 0.320 ;
        RECT 18.920 0.230 19.370 0.320 ;
        RECT 22.760 0.970 23.210 1.060 ;
        RECT 25.610 0.970 26.070 1.050 ;
        RECT 22.760 0.740 26.070 0.970 ;
        RECT 22.760 0.550 23.210 0.740 ;
        RECT 25.610 0.550 26.070 0.740 ;
        RECT 22.760 0.320 26.070 0.550 ;
        RECT 22.760 0.230 23.210 0.320 ;
        RECT 25.610 0.240 26.070 0.320 ;
        RECT 29.560 0.970 30.020 1.050 ;
        RECT 32.420 0.970 32.870 1.060 ;
        RECT 29.560 0.740 32.870 0.970 ;
        RECT 29.560 0.550 30.020 0.740 ;
        RECT 32.420 0.550 32.870 0.740 ;
        RECT 29.560 0.320 32.870 0.550 ;
        RECT 29.560 0.240 30.020 0.320 ;
        RECT 32.420 0.230 32.870 0.320 ;
        RECT 36.260 0.970 36.710 1.060 ;
        RECT 39.110 0.970 39.570 1.050 ;
        RECT 36.260 0.740 39.570 0.970 ;
        RECT 36.260 0.550 36.710 0.740 ;
        RECT 39.110 0.550 39.570 0.740 ;
        RECT 36.260 0.320 39.570 0.550 ;
        RECT 36.260 0.230 36.710 0.320 ;
        RECT 39.110 0.240 39.570 0.320 ;
        RECT 43.060 0.970 43.520 1.050 ;
        RECT 45.920 0.970 46.370 1.060 ;
        RECT 43.060 0.740 46.370 0.970 ;
        RECT 43.060 0.550 43.520 0.740 ;
        RECT 45.920 0.550 46.370 0.740 ;
        RECT 43.060 0.320 46.370 0.550 ;
        RECT 43.060 0.240 43.520 0.320 ;
        RECT 45.920 0.230 46.370 0.320 ;
        RECT 49.760 0.970 50.210 1.060 ;
        RECT 52.610 0.970 53.070 1.050 ;
        RECT 49.760 0.740 53.070 0.970 ;
        RECT 49.760 0.550 50.210 0.740 ;
        RECT 52.610 0.550 53.070 0.740 ;
        RECT 49.760 0.320 53.070 0.550 ;
        RECT 49.760 0.230 50.210 0.320 ;
        RECT 52.610 0.240 53.070 0.320 ;
        RECT 56.560 0.970 57.020 1.050 ;
        RECT 59.420 0.970 59.870 1.060 ;
        RECT 56.560 0.740 59.870 0.970 ;
        RECT 56.560 0.550 57.020 0.740 ;
        RECT 59.420 0.550 59.870 0.740 ;
        RECT 56.560 0.320 59.870 0.550 ;
        RECT 56.560 0.240 57.020 0.320 ;
        RECT 59.420 0.230 59.870 0.320 ;
        RECT 63.260 0.970 63.710 1.060 ;
        RECT 66.110 0.970 66.570 1.050 ;
        RECT 63.260 0.740 66.570 0.970 ;
        RECT 63.260 0.550 63.710 0.740 ;
        RECT 66.110 0.550 66.570 0.740 ;
        RECT 63.260 0.320 66.570 0.550 ;
        RECT 63.260 0.230 63.710 0.320 ;
        RECT 66.110 0.240 66.570 0.320 ;
        RECT 70.060 0.970 70.520 1.050 ;
        RECT 72.920 0.970 73.370 1.060 ;
        RECT 70.060 0.740 73.370 0.970 ;
        RECT 70.060 0.550 70.520 0.740 ;
        RECT 72.920 0.550 73.370 0.740 ;
        RECT 70.060 0.320 73.370 0.550 ;
        RECT 70.060 0.240 70.520 0.320 ;
        RECT 72.920 0.230 73.370 0.320 ;
        RECT 76.760 0.970 77.210 1.060 ;
        RECT 79.610 0.970 80.070 1.050 ;
        RECT 76.760 0.740 80.070 0.970 ;
        RECT 76.760 0.550 77.210 0.740 ;
        RECT 79.610 0.550 80.070 0.740 ;
        RECT 76.760 0.320 80.070 0.550 ;
        RECT 76.760 0.230 77.210 0.320 ;
        RECT 79.610 0.240 80.070 0.320 ;
        RECT 83.560 0.970 84.020 1.050 ;
        RECT 86.420 0.970 86.870 1.060 ;
        RECT 83.560 0.740 86.870 0.970 ;
        RECT 83.560 0.550 84.020 0.740 ;
        RECT 86.420 0.550 86.870 0.740 ;
        RECT 83.560 0.320 86.870 0.550 ;
        RECT 83.560 0.240 84.020 0.320 ;
        RECT 86.420 0.230 86.870 0.320 ;
        RECT 90.260 0.970 90.710 1.060 ;
        RECT 93.110 0.970 93.570 1.050 ;
        RECT 90.260 0.740 93.570 0.970 ;
        RECT 90.260 0.550 90.710 0.740 ;
        RECT 93.110 0.550 93.570 0.740 ;
        RECT 90.260 0.320 93.570 0.550 ;
        RECT 90.260 0.230 90.710 0.320 ;
        RECT 93.110 0.240 93.570 0.320 ;
        RECT 97.060 0.970 97.520 1.050 ;
        RECT 99.920 0.970 100.370 1.060 ;
        RECT 97.060 0.740 100.370 0.970 ;
        RECT 97.060 0.550 97.520 0.740 ;
        RECT 99.920 0.550 100.370 0.740 ;
        RECT 97.060 0.320 100.370 0.550 ;
        RECT 97.060 0.240 97.520 0.320 ;
        RECT 99.920 0.230 100.370 0.320 ;
        RECT 103.760 0.970 104.210 1.060 ;
        RECT 106.610 0.970 107.070 1.050 ;
        RECT 103.760 0.740 107.070 0.970 ;
        RECT 103.760 0.550 104.210 0.740 ;
        RECT 106.610 0.550 107.070 0.740 ;
        RECT 103.760 0.320 107.070 0.550 ;
        RECT 103.760 0.230 104.210 0.320 ;
        RECT 106.610 0.240 107.070 0.320 ;
        RECT 110.560 0.970 111.020 1.050 ;
        RECT 113.420 0.970 113.870 1.060 ;
        RECT 110.560 0.740 113.870 0.970 ;
        RECT 110.560 0.550 111.020 0.740 ;
        RECT 113.420 0.550 113.870 0.740 ;
        RECT 110.560 0.320 113.870 0.550 ;
        RECT 110.560 0.240 111.020 0.320 ;
        RECT 113.420 0.230 113.870 0.320 ;
        RECT 117.260 0.970 117.710 1.060 ;
        RECT 120.110 0.970 120.570 1.050 ;
        RECT 117.260 0.740 120.570 0.970 ;
        RECT 117.260 0.550 117.710 0.740 ;
        RECT 120.110 0.550 120.570 0.740 ;
        RECT 117.260 0.320 120.570 0.550 ;
        RECT 117.260 0.230 117.710 0.320 ;
        RECT 120.110 0.240 120.570 0.320 ;
        RECT 124.060 0.970 124.520 1.050 ;
        RECT 126.920 0.970 127.370 1.060 ;
        RECT 124.060 0.740 127.370 0.970 ;
        RECT 124.060 0.550 124.520 0.740 ;
        RECT 126.920 0.550 127.370 0.740 ;
        RECT 124.060 0.320 127.370 0.550 ;
        RECT 124.060 0.240 124.520 0.320 ;
        RECT 126.920 0.230 127.370 0.320 ;
        RECT 130.760 0.970 131.210 1.060 ;
        RECT 133.610 0.970 134.070 1.050 ;
        RECT 130.760 0.740 134.070 0.970 ;
        RECT 130.760 0.550 131.210 0.740 ;
        RECT 133.610 0.550 134.070 0.740 ;
        RECT 130.760 0.320 134.070 0.550 ;
        RECT 130.760 0.230 131.210 0.320 ;
        RECT 133.610 0.240 134.070 0.320 ;
        RECT 137.560 0.970 138.020 1.050 ;
        RECT 140.420 0.970 140.870 1.060 ;
        RECT 137.560 0.740 140.870 0.970 ;
        RECT 137.560 0.550 138.020 0.740 ;
        RECT 140.420 0.550 140.870 0.740 ;
        RECT 137.560 0.320 140.870 0.550 ;
        RECT 137.560 0.240 138.020 0.320 ;
        RECT 140.420 0.230 140.870 0.320 ;
        RECT 144.260 0.970 144.710 1.060 ;
        RECT 147.110 0.970 147.570 1.050 ;
        RECT 144.260 0.740 147.570 0.970 ;
        RECT 144.260 0.550 144.710 0.740 ;
        RECT 147.110 0.550 147.570 0.740 ;
        RECT 144.260 0.320 147.570 0.550 ;
        RECT 144.260 0.230 144.710 0.320 ;
        RECT 147.110 0.240 147.570 0.320 ;
        RECT 151.060 0.970 151.520 1.050 ;
        RECT 153.920 0.970 154.370 1.060 ;
        RECT 151.060 0.740 154.370 0.970 ;
        RECT 151.060 0.550 151.520 0.740 ;
        RECT 153.920 0.550 154.370 0.740 ;
        RECT 151.060 0.320 154.370 0.550 ;
        RECT 151.060 0.240 151.520 0.320 ;
        RECT 153.920 0.230 154.370 0.320 ;
        RECT 157.760 0.970 158.210 1.060 ;
        RECT 160.610 0.970 161.070 1.050 ;
        RECT 157.760 0.740 161.070 0.970 ;
        RECT 157.760 0.550 158.210 0.740 ;
        RECT 160.610 0.550 161.070 0.740 ;
        RECT 157.760 0.320 161.070 0.550 ;
        RECT 157.760 0.230 158.210 0.320 ;
        RECT 160.610 0.240 161.070 0.320 ;
        RECT 164.560 0.970 165.020 1.050 ;
        RECT 167.420 0.970 167.870 1.060 ;
        RECT 164.560 0.740 167.870 0.970 ;
        RECT 164.560 0.550 165.020 0.740 ;
        RECT 167.420 0.550 167.870 0.740 ;
        RECT 164.560 0.320 167.870 0.550 ;
        RECT 164.560 0.240 165.020 0.320 ;
        RECT 167.420 0.230 167.870 0.320 ;
        RECT 171.260 0.970 171.710 1.060 ;
        RECT 174.110 0.970 174.570 1.050 ;
        RECT 171.260 0.740 174.570 0.970 ;
        RECT 171.260 0.550 171.710 0.740 ;
        RECT 174.110 0.550 174.570 0.740 ;
        RECT 171.260 0.320 174.570 0.550 ;
        RECT 171.260 0.230 171.710 0.320 ;
        RECT 174.110 0.240 174.570 0.320 ;
        RECT 178.060 0.970 178.520 1.050 ;
        RECT 180.920 0.970 181.370 1.060 ;
        RECT 178.060 0.740 181.370 0.970 ;
        RECT 178.060 0.550 178.520 0.740 ;
        RECT 180.920 0.550 181.370 0.740 ;
        RECT 178.060 0.320 181.370 0.550 ;
        RECT 178.060 0.240 178.520 0.320 ;
        RECT 180.920 0.230 181.370 0.320 ;
        RECT 184.760 0.970 185.210 1.060 ;
        RECT 187.610 0.970 188.070 1.050 ;
        RECT 184.760 0.740 188.070 0.970 ;
        RECT 184.760 0.550 185.210 0.740 ;
        RECT 187.610 0.550 188.070 0.740 ;
        RECT 184.760 0.320 188.070 0.550 ;
        RECT 184.760 0.230 185.210 0.320 ;
        RECT 187.610 0.240 188.070 0.320 ;
        RECT 191.560 0.970 192.020 1.050 ;
        RECT 194.420 0.970 194.870 1.060 ;
        RECT 191.560 0.740 194.870 0.970 ;
        RECT 191.560 0.550 192.020 0.740 ;
        RECT 194.420 0.550 194.870 0.740 ;
        RECT 191.560 0.320 194.870 0.550 ;
        RECT 191.560 0.240 192.020 0.320 ;
        RECT 194.420 0.230 194.870 0.320 ;
        RECT 198.260 0.970 198.710 1.060 ;
        RECT 201.110 0.970 201.570 1.050 ;
        RECT 198.260 0.740 201.570 0.970 ;
        RECT 198.260 0.550 198.710 0.740 ;
        RECT 201.110 0.550 201.570 0.740 ;
        RECT 198.260 0.320 201.570 0.550 ;
        RECT 198.260 0.230 198.710 0.320 ;
        RECT 201.110 0.240 201.570 0.320 ;
        RECT 205.060 0.970 205.520 1.050 ;
        RECT 207.920 0.970 208.370 1.060 ;
        RECT 205.060 0.740 208.370 0.970 ;
        RECT 205.060 0.550 205.520 0.740 ;
        RECT 207.920 0.550 208.370 0.740 ;
        RECT 205.060 0.320 208.370 0.550 ;
        RECT 205.060 0.240 205.520 0.320 ;
        RECT 207.920 0.230 208.370 0.320 ;
        RECT 211.760 0.970 212.210 1.060 ;
        RECT 214.610 0.970 215.070 1.050 ;
        RECT 211.760 0.740 215.070 0.970 ;
        RECT 211.760 0.550 212.210 0.740 ;
        RECT 214.610 0.550 215.070 0.740 ;
        RECT 211.760 0.320 215.070 0.550 ;
        RECT 211.760 0.230 212.210 0.320 ;
        RECT 214.610 0.240 215.070 0.320 ;
        RECT 9.260 -2.640 9.710 -2.550 ;
        RECT 12.110 -2.640 12.570 -2.560 ;
        RECT 9.260 -2.870 12.570 -2.640 ;
        RECT 9.260 -3.060 9.710 -2.870 ;
        RECT 12.110 -3.060 12.570 -2.870 ;
        RECT 9.260 -3.290 12.570 -3.060 ;
        RECT 9.260 -3.380 9.710 -3.290 ;
        RECT 12.110 -3.370 12.570 -3.290 ;
        RECT 16.060 -2.640 16.520 -2.560 ;
        RECT 18.920 -2.640 19.370 -2.550 ;
        RECT 16.060 -2.870 19.370 -2.640 ;
        RECT 16.060 -3.060 16.520 -2.870 ;
        RECT 18.920 -3.060 19.370 -2.870 ;
        RECT 16.060 -3.290 19.370 -3.060 ;
        RECT 16.060 -3.370 16.520 -3.290 ;
        RECT 18.920 -3.380 19.370 -3.290 ;
        RECT 22.760 -2.640 23.210 -2.550 ;
        RECT 25.610 -2.640 26.070 -2.560 ;
        RECT 22.760 -2.870 26.070 -2.640 ;
        RECT 22.760 -3.060 23.210 -2.870 ;
        RECT 25.610 -3.060 26.070 -2.870 ;
        RECT 22.760 -3.290 26.070 -3.060 ;
        RECT 22.760 -3.380 23.210 -3.290 ;
        RECT 25.610 -3.370 26.070 -3.290 ;
        RECT 29.560 -2.640 30.020 -2.560 ;
        RECT 32.420 -2.640 32.870 -2.550 ;
        RECT 29.560 -2.870 32.870 -2.640 ;
        RECT 29.560 -3.060 30.020 -2.870 ;
        RECT 32.420 -3.060 32.870 -2.870 ;
        RECT 29.560 -3.290 32.870 -3.060 ;
        RECT 29.560 -3.370 30.020 -3.290 ;
        RECT 32.420 -3.380 32.870 -3.290 ;
        RECT 36.260 -2.640 36.710 -2.550 ;
        RECT 39.110 -2.640 39.570 -2.560 ;
        RECT 36.260 -2.870 39.570 -2.640 ;
        RECT 36.260 -3.060 36.710 -2.870 ;
        RECT 39.110 -3.060 39.570 -2.870 ;
        RECT 36.260 -3.290 39.570 -3.060 ;
        RECT 36.260 -3.380 36.710 -3.290 ;
        RECT 39.110 -3.370 39.570 -3.290 ;
        RECT 43.060 -2.640 43.520 -2.560 ;
        RECT 45.920 -2.640 46.370 -2.550 ;
        RECT 43.060 -2.870 46.370 -2.640 ;
        RECT 43.060 -3.060 43.520 -2.870 ;
        RECT 45.920 -3.060 46.370 -2.870 ;
        RECT 43.060 -3.290 46.370 -3.060 ;
        RECT 43.060 -3.370 43.520 -3.290 ;
        RECT 45.920 -3.380 46.370 -3.290 ;
        RECT 49.760 -2.640 50.210 -2.550 ;
        RECT 52.610 -2.640 53.070 -2.560 ;
        RECT 49.760 -2.870 53.070 -2.640 ;
        RECT 49.760 -3.060 50.210 -2.870 ;
        RECT 52.610 -3.060 53.070 -2.870 ;
        RECT 49.760 -3.290 53.070 -3.060 ;
        RECT 49.760 -3.380 50.210 -3.290 ;
        RECT 52.610 -3.370 53.070 -3.290 ;
        RECT 56.560 -2.640 57.020 -2.560 ;
        RECT 59.420 -2.640 59.870 -2.550 ;
        RECT 56.560 -2.870 59.870 -2.640 ;
        RECT 56.560 -3.060 57.020 -2.870 ;
        RECT 59.420 -3.060 59.870 -2.870 ;
        RECT 56.560 -3.290 59.870 -3.060 ;
        RECT 56.560 -3.370 57.020 -3.290 ;
        RECT 59.420 -3.380 59.870 -3.290 ;
        RECT 63.260 -2.640 63.710 -2.550 ;
        RECT 66.110 -2.640 66.570 -2.560 ;
        RECT 63.260 -2.870 66.570 -2.640 ;
        RECT 63.260 -3.060 63.710 -2.870 ;
        RECT 66.110 -3.060 66.570 -2.870 ;
        RECT 63.260 -3.290 66.570 -3.060 ;
        RECT 63.260 -3.380 63.710 -3.290 ;
        RECT 66.110 -3.370 66.570 -3.290 ;
        RECT 70.060 -2.640 70.520 -2.560 ;
        RECT 72.920 -2.640 73.370 -2.550 ;
        RECT 70.060 -2.870 73.370 -2.640 ;
        RECT 70.060 -3.060 70.520 -2.870 ;
        RECT 72.920 -3.060 73.370 -2.870 ;
        RECT 70.060 -3.290 73.370 -3.060 ;
        RECT 70.060 -3.370 70.520 -3.290 ;
        RECT 72.920 -3.380 73.370 -3.290 ;
        RECT 76.760 -2.640 77.210 -2.550 ;
        RECT 79.610 -2.640 80.070 -2.560 ;
        RECT 76.760 -2.870 80.070 -2.640 ;
        RECT 76.760 -3.060 77.210 -2.870 ;
        RECT 79.610 -3.060 80.070 -2.870 ;
        RECT 76.760 -3.290 80.070 -3.060 ;
        RECT 76.760 -3.380 77.210 -3.290 ;
        RECT 79.610 -3.370 80.070 -3.290 ;
        RECT 83.560 -2.640 84.020 -2.560 ;
        RECT 86.420 -2.640 86.870 -2.550 ;
        RECT 83.560 -2.870 86.870 -2.640 ;
        RECT 83.560 -3.060 84.020 -2.870 ;
        RECT 86.420 -3.060 86.870 -2.870 ;
        RECT 83.560 -3.290 86.870 -3.060 ;
        RECT 83.560 -3.370 84.020 -3.290 ;
        RECT 86.420 -3.380 86.870 -3.290 ;
        RECT 90.260 -2.640 90.710 -2.550 ;
        RECT 93.110 -2.640 93.570 -2.560 ;
        RECT 90.260 -2.870 93.570 -2.640 ;
        RECT 90.260 -3.060 90.710 -2.870 ;
        RECT 93.110 -3.060 93.570 -2.870 ;
        RECT 90.260 -3.290 93.570 -3.060 ;
        RECT 90.260 -3.380 90.710 -3.290 ;
        RECT 93.110 -3.370 93.570 -3.290 ;
        RECT 97.060 -2.640 97.520 -2.560 ;
        RECT 99.920 -2.640 100.370 -2.550 ;
        RECT 97.060 -2.870 100.370 -2.640 ;
        RECT 97.060 -3.060 97.520 -2.870 ;
        RECT 99.920 -3.060 100.370 -2.870 ;
        RECT 97.060 -3.290 100.370 -3.060 ;
        RECT 97.060 -3.370 97.520 -3.290 ;
        RECT 99.920 -3.380 100.370 -3.290 ;
        RECT 103.760 -2.640 104.210 -2.550 ;
        RECT 106.610 -2.640 107.070 -2.560 ;
        RECT 103.760 -2.870 107.070 -2.640 ;
        RECT 103.760 -3.060 104.210 -2.870 ;
        RECT 106.610 -3.060 107.070 -2.870 ;
        RECT 103.760 -3.290 107.070 -3.060 ;
        RECT 103.760 -3.380 104.210 -3.290 ;
        RECT 106.610 -3.370 107.070 -3.290 ;
        RECT 110.560 -2.640 111.020 -2.560 ;
        RECT 113.420 -2.640 113.870 -2.550 ;
        RECT 110.560 -2.870 113.870 -2.640 ;
        RECT 110.560 -3.060 111.020 -2.870 ;
        RECT 113.420 -3.060 113.870 -2.870 ;
        RECT 110.560 -3.290 113.870 -3.060 ;
        RECT 110.560 -3.370 111.020 -3.290 ;
        RECT 113.420 -3.380 113.870 -3.290 ;
        RECT 117.260 -2.640 117.710 -2.550 ;
        RECT 120.110 -2.640 120.570 -2.560 ;
        RECT 117.260 -2.870 120.570 -2.640 ;
        RECT 117.260 -3.060 117.710 -2.870 ;
        RECT 120.110 -3.060 120.570 -2.870 ;
        RECT 117.260 -3.290 120.570 -3.060 ;
        RECT 117.260 -3.380 117.710 -3.290 ;
        RECT 120.110 -3.370 120.570 -3.290 ;
        RECT 124.060 -2.640 124.520 -2.560 ;
        RECT 126.920 -2.640 127.370 -2.550 ;
        RECT 124.060 -2.870 127.370 -2.640 ;
        RECT 124.060 -3.060 124.520 -2.870 ;
        RECT 126.920 -3.060 127.370 -2.870 ;
        RECT 124.060 -3.290 127.370 -3.060 ;
        RECT 124.060 -3.370 124.520 -3.290 ;
        RECT 126.920 -3.380 127.370 -3.290 ;
        RECT 130.760 -2.640 131.210 -2.550 ;
        RECT 133.610 -2.640 134.070 -2.560 ;
        RECT 130.760 -2.870 134.070 -2.640 ;
        RECT 130.760 -3.060 131.210 -2.870 ;
        RECT 133.610 -3.060 134.070 -2.870 ;
        RECT 130.760 -3.290 134.070 -3.060 ;
        RECT 130.760 -3.380 131.210 -3.290 ;
        RECT 133.610 -3.370 134.070 -3.290 ;
        RECT 137.560 -2.640 138.020 -2.560 ;
        RECT 140.420 -2.640 140.870 -2.550 ;
        RECT 137.560 -2.870 140.870 -2.640 ;
        RECT 137.560 -3.060 138.020 -2.870 ;
        RECT 140.420 -3.060 140.870 -2.870 ;
        RECT 137.560 -3.290 140.870 -3.060 ;
        RECT 137.560 -3.370 138.020 -3.290 ;
        RECT 140.420 -3.380 140.870 -3.290 ;
        RECT 144.260 -2.640 144.710 -2.550 ;
        RECT 147.110 -2.640 147.570 -2.560 ;
        RECT 144.260 -2.870 147.570 -2.640 ;
        RECT 144.260 -3.060 144.710 -2.870 ;
        RECT 147.110 -3.060 147.570 -2.870 ;
        RECT 144.260 -3.290 147.570 -3.060 ;
        RECT 144.260 -3.380 144.710 -3.290 ;
        RECT 147.110 -3.370 147.570 -3.290 ;
        RECT 151.060 -2.640 151.520 -2.560 ;
        RECT 153.920 -2.640 154.370 -2.550 ;
        RECT 151.060 -2.870 154.370 -2.640 ;
        RECT 151.060 -3.060 151.520 -2.870 ;
        RECT 153.920 -3.060 154.370 -2.870 ;
        RECT 151.060 -3.290 154.370 -3.060 ;
        RECT 151.060 -3.370 151.520 -3.290 ;
        RECT 153.920 -3.380 154.370 -3.290 ;
        RECT 157.760 -2.640 158.210 -2.550 ;
        RECT 160.610 -2.640 161.070 -2.560 ;
        RECT 157.760 -2.870 161.070 -2.640 ;
        RECT 157.760 -3.060 158.210 -2.870 ;
        RECT 160.610 -3.060 161.070 -2.870 ;
        RECT 157.760 -3.290 161.070 -3.060 ;
        RECT 157.760 -3.380 158.210 -3.290 ;
        RECT 160.610 -3.370 161.070 -3.290 ;
        RECT 164.560 -2.640 165.020 -2.560 ;
        RECT 167.420 -2.640 167.870 -2.550 ;
        RECT 164.560 -2.870 167.870 -2.640 ;
        RECT 164.560 -3.060 165.020 -2.870 ;
        RECT 167.420 -3.060 167.870 -2.870 ;
        RECT 164.560 -3.290 167.870 -3.060 ;
        RECT 164.560 -3.370 165.020 -3.290 ;
        RECT 167.420 -3.380 167.870 -3.290 ;
        RECT 171.260 -2.640 171.710 -2.550 ;
        RECT 174.110 -2.640 174.570 -2.560 ;
        RECT 171.260 -2.870 174.570 -2.640 ;
        RECT 171.260 -3.060 171.710 -2.870 ;
        RECT 174.110 -3.060 174.570 -2.870 ;
        RECT 171.260 -3.290 174.570 -3.060 ;
        RECT 171.260 -3.380 171.710 -3.290 ;
        RECT 174.110 -3.370 174.570 -3.290 ;
        RECT 178.060 -2.640 178.520 -2.560 ;
        RECT 180.920 -2.640 181.370 -2.550 ;
        RECT 178.060 -2.870 181.370 -2.640 ;
        RECT 178.060 -3.060 178.520 -2.870 ;
        RECT 180.920 -3.060 181.370 -2.870 ;
        RECT 178.060 -3.290 181.370 -3.060 ;
        RECT 178.060 -3.370 178.520 -3.290 ;
        RECT 180.920 -3.380 181.370 -3.290 ;
        RECT 184.760 -2.640 185.210 -2.550 ;
        RECT 187.610 -2.640 188.070 -2.560 ;
        RECT 184.760 -2.870 188.070 -2.640 ;
        RECT 184.760 -3.060 185.210 -2.870 ;
        RECT 187.610 -3.060 188.070 -2.870 ;
        RECT 184.760 -3.290 188.070 -3.060 ;
        RECT 184.760 -3.380 185.210 -3.290 ;
        RECT 187.610 -3.370 188.070 -3.290 ;
        RECT 191.560 -2.640 192.020 -2.560 ;
        RECT 194.420 -2.640 194.870 -2.550 ;
        RECT 191.560 -2.870 194.870 -2.640 ;
        RECT 191.560 -3.060 192.020 -2.870 ;
        RECT 194.420 -3.060 194.870 -2.870 ;
        RECT 191.560 -3.290 194.870 -3.060 ;
        RECT 191.560 -3.370 192.020 -3.290 ;
        RECT 194.420 -3.380 194.870 -3.290 ;
        RECT 198.260 -2.640 198.710 -2.550 ;
        RECT 201.110 -2.640 201.570 -2.560 ;
        RECT 198.260 -2.870 201.570 -2.640 ;
        RECT 198.260 -3.060 198.710 -2.870 ;
        RECT 201.110 -3.060 201.570 -2.870 ;
        RECT 198.260 -3.290 201.570 -3.060 ;
        RECT 198.260 -3.380 198.710 -3.290 ;
        RECT 201.110 -3.370 201.570 -3.290 ;
        RECT 205.060 -2.640 205.520 -2.560 ;
        RECT 207.920 -2.640 208.370 -2.550 ;
        RECT 205.060 -2.870 208.370 -2.640 ;
        RECT 205.060 -3.060 205.520 -2.870 ;
        RECT 207.920 -3.060 208.370 -2.870 ;
        RECT 205.060 -3.290 208.370 -3.060 ;
        RECT 205.060 -3.370 205.520 -3.290 ;
        RECT 207.920 -3.380 208.370 -3.290 ;
        RECT 211.760 -2.640 212.210 -2.550 ;
        RECT 214.610 -2.640 215.070 -2.560 ;
        RECT 211.760 -2.870 215.070 -2.640 ;
        RECT 211.760 -3.060 212.210 -2.870 ;
        RECT 214.610 -3.060 215.070 -2.870 ;
        RECT 211.760 -3.290 215.070 -3.060 ;
        RECT 211.760 -3.380 212.210 -3.290 ;
        RECT 214.610 -3.370 215.070 -3.290 ;
        RECT 9.260 -6.250 9.710 -6.160 ;
        RECT 12.110 -6.250 12.570 -6.170 ;
        RECT 9.260 -6.480 12.570 -6.250 ;
        RECT 9.260 -6.670 9.710 -6.480 ;
        RECT 12.110 -6.670 12.570 -6.480 ;
        RECT 9.260 -6.900 12.570 -6.670 ;
        RECT 9.260 -6.990 9.710 -6.900 ;
        RECT 12.110 -6.980 12.570 -6.900 ;
        RECT 16.060 -6.250 16.520 -6.170 ;
        RECT 18.920 -6.250 19.370 -6.160 ;
        RECT 16.060 -6.480 19.370 -6.250 ;
        RECT 16.060 -6.670 16.520 -6.480 ;
        RECT 18.920 -6.670 19.370 -6.480 ;
        RECT 16.060 -6.900 19.370 -6.670 ;
        RECT 16.060 -6.980 16.520 -6.900 ;
        RECT 18.920 -6.990 19.370 -6.900 ;
        RECT 22.760 -6.250 23.210 -6.160 ;
        RECT 25.610 -6.250 26.070 -6.170 ;
        RECT 22.760 -6.480 26.070 -6.250 ;
        RECT 22.760 -6.670 23.210 -6.480 ;
        RECT 25.610 -6.670 26.070 -6.480 ;
        RECT 22.760 -6.900 26.070 -6.670 ;
        RECT 22.760 -6.990 23.210 -6.900 ;
        RECT 25.610 -6.980 26.070 -6.900 ;
        RECT 29.560 -6.250 30.020 -6.170 ;
        RECT 32.420 -6.250 32.870 -6.160 ;
        RECT 29.560 -6.480 32.870 -6.250 ;
        RECT 29.560 -6.670 30.020 -6.480 ;
        RECT 32.420 -6.670 32.870 -6.480 ;
        RECT 29.560 -6.900 32.870 -6.670 ;
        RECT 29.560 -6.980 30.020 -6.900 ;
        RECT 32.420 -6.990 32.870 -6.900 ;
        RECT 36.260 -6.250 36.710 -6.160 ;
        RECT 39.110 -6.250 39.570 -6.170 ;
        RECT 36.260 -6.480 39.570 -6.250 ;
        RECT 36.260 -6.670 36.710 -6.480 ;
        RECT 39.110 -6.670 39.570 -6.480 ;
        RECT 36.260 -6.900 39.570 -6.670 ;
        RECT 36.260 -6.990 36.710 -6.900 ;
        RECT 39.110 -6.980 39.570 -6.900 ;
        RECT 43.060 -6.250 43.520 -6.170 ;
        RECT 45.920 -6.250 46.370 -6.160 ;
        RECT 43.060 -6.480 46.370 -6.250 ;
        RECT 43.060 -6.670 43.520 -6.480 ;
        RECT 45.920 -6.670 46.370 -6.480 ;
        RECT 43.060 -6.900 46.370 -6.670 ;
        RECT 43.060 -6.980 43.520 -6.900 ;
        RECT 45.920 -6.990 46.370 -6.900 ;
        RECT 49.760 -6.250 50.210 -6.160 ;
        RECT 52.610 -6.250 53.070 -6.170 ;
        RECT 49.760 -6.480 53.070 -6.250 ;
        RECT 49.760 -6.670 50.210 -6.480 ;
        RECT 52.610 -6.670 53.070 -6.480 ;
        RECT 49.760 -6.900 53.070 -6.670 ;
        RECT 49.760 -6.990 50.210 -6.900 ;
        RECT 52.610 -6.980 53.070 -6.900 ;
        RECT 56.560 -6.250 57.020 -6.170 ;
        RECT 59.420 -6.250 59.870 -6.160 ;
        RECT 56.560 -6.480 59.870 -6.250 ;
        RECT 56.560 -6.670 57.020 -6.480 ;
        RECT 59.420 -6.670 59.870 -6.480 ;
        RECT 56.560 -6.900 59.870 -6.670 ;
        RECT 56.560 -6.980 57.020 -6.900 ;
        RECT 59.420 -6.990 59.870 -6.900 ;
        RECT 63.260 -6.250 63.710 -6.160 ;
        RECT 66.110 -6.250 66.570 -6.170 ;
        RECT 63.260 -6.480 66.570 -6.250 ;
        RECT 63.260 -6.670 63.710 -6.480 ;
        RECT 66.110 -6.670 66.570 -6.480 ;
        RECT 63.260 -6.900 66.570 -6.670 ;
        RECT 63.260 -6.990 63.710 -6.900 ;
        RECT 66.110 -6.980 66.570 -6.900 ;
        RECT 70.060 -6.250 70.520 -6.170 ;
        RECT 72.920 -6.250 73.370 -6.160 ;
        RECT 70.060 -6.480 73.370 -6.250 ;
        RECT 70.060 -6.670 70.520 -6.480 ;
        RECT 72.920 -6.670 73.370 -6.480 ;
        RECT 70.060 -6.900 73.370 -6.670 ;
        RECT 70.060 -6.980 70.520 -6.900 ;
        RECT 72.920 -6.990 73.370 -6.900 ;
        RECT 76.760 -6.250 77.210 -6.160 ;
        RECT 79.610 -6.250 80.070 -6.170 ;
        RECT 76.760 -6.480 80.070 -6.250 ;
        RECT 76.760 -6.670 77.210 -6.480 ;
        RECT 79.610 -6.670 80.070 -6.480 ;
        RECT 76.760 -6.900 80.070 -6.670 ;
        RECT 76.760 -6.990 77.210 -6.900 ;
        RECT 79.610 -6.980 80.070 -6.900 ;
        RECT 83.560 -6.250 84.020 -6.170 ;
        RECT 86.420 -6.250 86.870 -6.160 ;
        RECT 83.560 -6.480 86.870 -6.250 ;
        RECT 83.560 -6.670 84.020 -6.480 ;
        RECT 86.420 -6.670 86.870 -6.480 ;
        RECT 83.560 -6.900 86.870 -6.670 ;
        RECT 83.560 -6.980 84.020 -6.900 ;
        RECT 86.420 -6.990 86.870 -6.900 ;
        RECT 90.260 -6.250 90.710 -6.160 ;
        RECT 93.110 -6.250 93.570 -6.170 ;
        RECT 90.260 -6.480 93.570 -6.250 ;
        RECT 90.260 -6.670 90.710 -6.480 ;
        RECT 93.110 -6.670 93.570 -6.480 ;
        RECT 90.260 -6.900 93.570 -6.670 ;
        RECT 90.260 -6.990 90.710 -6.900 ;
        RECT 93.110 -6.980 93.570 -6.900 ;
        RECT 97.060 -6.250 97.520 -6.170 ;
        RECT 99.920 -6.250 100.370 -6.160 ;
        RECT 97.060 -6.480 100.370 -6.250 ;
        RECT 97.060 -6.670 97.520 -6.480 ;
        RECT 99.920 -6.670 100.370 -6.480 ;
        RECT 97.060 -6.900 100.370 -6.670 ;
        RECT 97.060 -6.980 97.520 -6.900 ;
        RECT 99.920 -6.990 100.370 -6.900 ;
        RECT 103.760 -6.250 104.210 -6.160 ;
        RECT 106.610 -6.250 107.070 -6.170 ;
        RECT 103.760 -6.480 107.070 -6.250 ;
        RECT 103.760 -6.670 104.210 -6.480 ;
        RECT 106.610 -6.670 107.070 -6.480 ;
        RECT 103.760 -6.900 107.070 -6.670 ;
        RECT 103.760 -6.990 104.210 -6.900 ;
        RECT 106.610 -6.980 107.070 -6.900 ;
        RECT 110.560 -6.250 111.020 -6.170 ;
        RECT 113.420 -6.250 113.870 -6.160 ;
        RECT 110.560 -6.480 113.870 -6.250 ;
        RECT 110.560 -6.670 111.020 -6.480 ;
        RECT 113.420 -6.670 113.870 -6.480 ;
        RECT 110.560 -6.900 113.870 -6.670 ;
        RECT 110.560 -6.980 111.020 -6.900 ;
        RECT 113.420 -6.990 113.870 -6.900 ;
        RECT 117.260 -6.250 117.710 -6.160 ;
        RECT 120.110 -6.250 120.570 -6.170 ;
        RECT 117.260 -6.480 120.570 -6.250 ;
        RECT 117.260 -6.670 117.710 -6.480 ;
        RECT 120.110 -6.670 120.570 -6.480 ;
        RECT 117.260 -6.900 120.570 -6.670 ;
        RECT 117.260 -6.990 117.710 -6.900 ;
        RECT 120.110 -6.980 120.570 -6.900 ;
        RECT 124.060 -6.250 124.520 -6.170 ;
        RECT 126.920 -6.250 127.370 -6.160 ;
        RECT 124.060 -6.480 127.370 -6.250 ;
        RECT 124.060 -6.670 124.520 -6.480 ;
        RECT 126.920 -6.670 127.370 -6.480 ;
        RECT 124.060 -6.900 127.370 -6.670 ;
        RECT 124.060 -6.980 124.520 -6.900 ;
        RECT 126.920 -6.990 127.370 -6.900 ;
        RECT 130.760 -6.250 131.210 -6.160 ;
        RECT 133.610 -6.250 134.070 -6.170 ;
        RECT 130.760 -6.480 134.070 -6.250 ;
        RECT 130.760 -6.670 131.210 -6.480 ;
        RECT 133.610 -6.670 134.070 -6.480 ;
        RECT 130.760 -6.900 134.070 -6.670 ;
        RECT 130.760 -6.990 131.210 -6.900 ;
        RECT 133.610 -6.980 134.070 -6.900 ;
        RECT 137.560 -6.250 138.020 -6.170 ;
        RECT 140.420 -6.250 140.870 -6.160 ;
        RECT 137.560 -6.480 140.870 -6.250 ;
        RECT 137.560 -6.670 138.020 -6.480 ;
        RECT 140.420 -6.670 140.870 -6.480 ;
        RECT 137.560 -6.900 140.870 -6.670 ;
        RECT 137.560 -6.980 138.020 -6.900 ;
        RECT 140.420 -6.990 140.870 -6.900 ;
        RECT 144.260 -6.250 144.710 -6.160 ;
        RECT 147.110 -6.250 147.570 -6.170 ;
        RECT 144.260 -6.480 147.570 -6.250 ;
        RECT 144.260 -6.670 144.710 -6.480 ;
        RECT 147.110 -6.670 147.570 -6.480 ;
        RECT 144.260 -6.900 147.570 -6.670 ;
        RECT 144.260 -6.990 144.710 -6.900 ;
        RECT 147.110 -6.980 147.570 -6.900 ;
        RECT 151.060 -6.250 151.520 -6.170 ;
        RECT 153.920 -6.250 154.370 -6.160 ;
        RECT 151.060 -6.480 154.370 -6.250 ;
        RECT 151.060 -6.670 151.520 -6.480 ;
        RECT 153.920 -6.670 154.370 -6.480 ;
        RECT 151.060 -6.900 154.370 -6.670 ;
        RECT 151.060 -6.980 151.520 -6.900 ;
        RECT 153.920 -6.990 154.370 -6.900 ;
        RECT 157.760 -6.250 158.210 -6.160 ;
        RECT 160.610 -6.250 161.070 -6.170 ;
        RECT 157.760 -6.480 161.070 -6.250 ;
        RECT 157.760 -6.670 158.210 -6.480 ;
        RECT 160.610 -6.670 161.070 -6.480 ;
        RECT 157.760 -6.900 161.070 -6.670 ;
        RECT 157.760 -6.990 158.210 -6.900 ;
        RECT 160.610 -6.980 161.070 -6.900 ;
        RECT 164.560 -6.250 165.020 -6.170 ;
        RECT 167.420 -6.250 167.870 -6.160 ;
        RECT 164.560 -6.480 167.870 -6.250 ;
        RECT 164.560 -6.670 165.020 -6.480 ;
        RECT 167.420 -6.670 167.870 -6.480 ;
        RECT 164.560 -6.900 167.870 -6.670 ;
        RECT 164.560 -6.980 165.020 -6.900 ;
        RECT 167.420 -6.990 167.870 -6.900 ;
        RECT 171.260 -6.250 171.710 -6.160 ;
        RECT 174.110 -6.250 174.570 -6.170 ;
        RECT 171.260 -6.480 174.570 -6.250 ;
        RECT 171.260 -6.670 171.710 -6.480 ;
        RECT 174.110 -6.670 174.570 -6.480 ;
        RECT 171.260 -6.900 174.570 -6.670 ;
        RECT 171.260 -6.990 171.710 -6.900 ;
        RECT 174.110 -6.980 174.570 -6.900 ;
        RECT 178.060 -6.250 178.520 -6.170 ;
        RECT 180.920 -6.250 181.370 -6.160 ;
        RECT 178.060 -6.480 181.370 -6.250 ;
        RECT 178.060 -6.670 178.520 -6.480 ;
        RECT 180.920 -6.670 181.370 -6.480 ;
        RECT 178.060 -6.900 181.370 -6.670 ;
        RECT 178.060 -6.980 178.520 -6.900 ;
        RECT 180.920 -6.990 181.370 -6.900 ;
        RECT 184.760 -6.250 185.210 -6.160 ;
        RECT 187.610 -6.250 188.070 -6.170 ;
        RECT 184.760 -6.480 188.070 -6.250 ;
        RECT 184.760 -6.670 185.210 -6.480 ;
        RECT 187.610 -6.670 188.070 -6.480 ;
        RECT 184.760 -6.900 188.070 -6.670 ;
        RECT 184.760 -6.990 185.210 -6.900 ;
        RECT 187.610 -6.980 188.070 -6.900 ;
        RECT 191.560 -6.250 192.020 -6.170 ;
        RECT 194.420 -6.250 194.870 -6.160 ;
        RECT 191.560 -6.480 194.870 -6.250 ;
        RECT 191.560 -6.670 192.020 -6.480 ;
        RECT 194.420 -6.670 194.870 -6.480 ;
        RECT 191.560 -6.900 194.870 -6.670 ;
        RECT 191.560 -6.980 192.020 -6.900 ;
        RECT 194.420 -6.990 194.870 -6.900 ;
        RECT 198.260 -6.250 198.710 -6.160 ;
        RECT 201.110 -6.250 201.570 -6.170 ;
        RECT 198.260 -6.480 201.570 -6.250 ;
        RECT 198.260 -6.670 198.710 -6.480 ;
        RECT 201.110 -6.670 201.570 -6.480 ;
        RECT 198.260 -6.900 201.570 -6.670 ;
        RECT 198.260 -6.990 198.710 -6.900 ;
        RECT 201.110 -6.980 201.570 -6.900 ;
        RECT 205.060 -6.250 205.520 -6.170 ;
        RECT 207.920 -6.250 208.370 -6.160 ;
        RECT 205.060 -6.480 208.370 -6.250 ;
        RECT 205.060 -6.670 205.520 -6.480 ;
        RECT 207.920 -6.670 208.370 -6.480 ;
        RECT 205.060 -6.900 208.370 -6.670 ;
        RECT 205.060 -6.980 205.520 -6.900 ;
        RECT 207.920 -6.990 208.370 -6.900 ;
        RECT 211.760 -6.250 212.210 -6.160 ;
        RECT 214.610 -6.250 215.070 -6.170 ;
        RECT 211.760 -6.480 215.070 -6.250 ;
        RECT 211.760 -6.670 212.210 -6.480 ;
        RECT 214.610 -6.670 215.070 -6.480 ;
        RECT 211.760 -6.900 215.070 -6.670 ;
        RECT 211.760 -6.990 212.210 -6.900 ;
        RECT 214.610 -6.980 215.070 -6.900 ;
        RECT 9.260 -9.860 9.710 -9.770 ;
        RECT 12.110 -9.860 12.570 -9.780 ;
        RECT 9.260 -10.090 12.570 -9.860 ;
        RECT 9.260 -10.280 9.710 -10.090 ;
        RECT 12.110 -10.280 12.570 -10.090 ;
        RECT 9.260 -10.510 12.570 -10.280 ;
        RECT 9.260 -10.600 9.710 -10.510 ;
        RECT 12.110 -10.590 12.570 -10.510 ;
        RECT 16.060 -9.860 16.520 -9.780 ;
        RECT 18.920 -9.860 19.370 -9.770 ;
        RECT 16.060 -10.090 19.370 -9.860 ;
        RECT 16.060 -10.280 16.520 -10.090 ;
        RECT 18.920 -10.280 19.370 -10.090 ;
        RECT 16.060 -10.510 19.370 -10.280 ;
        RECT 16.060 -10.590 16.520 -10.510 ;
        RECT 18.920 -10.600 19.370 -10.510 ;
        RECT 22.760 -9.860 23.210 -9.770 ;
        RECT 25.610 -9.860 26.070 -9.780 ;
        RECT 22.760 -10.090 26.070 -9.860 ;
        RECT 22.760 -10.280 23.210 -10.090 ;
        RECT 25.610 -10.280 26.070 -10.090 ;
        RECT 22.760 -10.510 26.070 -10.280 ;
        RECT 22.760 -10.600 23.210 -10.510 ;
        RECT 25.610 -10.590 26.070 -10.510 ;
        RECT 29.560 -9.860 30.020 -9.780 ;
        RECT 32.420 -9.860 32.870 -9.770 ;
        RECT 29.560 -10.090 32.870 -9.860 ;
        RECT 29.560 -10.280 30.020 -10.090 ;
        RECT 32.420 -10.280 32.870 -10.090 ;
        RECT 29.560 -10.510 32.870 -10.280 ;
        RECT 29.560 -10.590 30.020 -10.510 ;
        RECT 32.420 -10.600 32.870 -10.510 ;
        RECT 36.260 -9.860 36.710 -9.770 ;
        RECT 39.110 -9.860 39.570 -9.780 ;
        RECT 36.260 -10.090 39.570 -9.860 ;
        RECT 36.260 -10.280 36.710 -10.090 ;
        RECT 39.110 -10.280 39.570 -10.090 ;
        RECT 36.260 -10.510 39.570 -10.280 ;
        RECT 36.260 -10.600 36.710 -10.510 ;
        RECT 39.110 -10.590 39.570 -10.510 ;
        RECT 43.060 -9.860 43.520 -9.780 ;
        RECT 45.920 -9.860 46.370 -9.770 ;
        RECT 43.060 -10.090 46.370 -9.860 ;
        RECT 43.060 -10.280 43.520 -10.090 ;
        RECT 45.920 -10.280 46.370 -10.090 ;
        RECT 43.060 -10.510 46.370 -10.280 ;
        RECT 43.060 -10.590 43.520 -10.510 ;
        RECT 45.920 -10.600 46.370 -10.510 ;
        RECT 49.760 -9.860 50.210 -9.770 ;
        RECT 52.610 -9.860 53.070 -9.780 ;
        RECT 49.760 -10.090 53.070 -9.860 ;
        RECT 49.760 -10.280 50.210 -10.090 ;
        RECT 52.610 -10.280 53.070 -10.090 ;
        RECT 49.760 -10.510 53.070 -10.280 ;
        RECT 49.760 -10.600 50.210 -10.510 ;
        RECT 52.610 -10.590 53.070 -10.510 ;
        RECT 56.560 -9.860 57.020 -9.780 ;
        RECT 59.420 -9.860 59.870 -9.770 ;
        RECT 56.560 -10.090 59.870 -9.860 ;
        RECT 56.560 -10.280 57.020 -10.090 ;
        RECT 59.420 -10.280 59.870 -10.090 ;
        RECT 56.560 -10.510 59.870 -10.280 ;
        RECT 56.560 -10.590 57.020 -10.510 ;
        RECT 59.420 -10.600 59.870 -10.510 ;
        RECT 63.260 -9.860 63.710 -9.770 ;
        RECT 66.110 -9.860 66.570 -9.780 ;
        RECT 63.260 -10.090 66.570 -9.860 ;
        RECT 63.260 -10.280 63.710 -10.090 ;
        RECT 66.110 -10.280 66.570 -10.090 ;
        RECT 63.260 -10.510 66.570 -10.280 ;
        RECT 63.260 -10.600 63.710 -10.510 ;
        RECT 66.110 -10.590 66.570 -10.510 ;
        RECT 70.060 -9.860 70.520 -9.780 ;
        RECT 72.920 -9.860 73.370 -9.770 ;
        RECT 70.060 -10.090 73.370 -9.860 ;
        RECT 70.060 -10.280 70.520 -10.090 ;
        RECT 72.920 -10.280 73.370 -10.090 ;
        RECT 70.060 -10.510 73.370 -10.280 ;
        RECT 70.060 -10.590 70.520 -10.510 ;
        RECT 72.920 -10.600 73.370 -10.510 ;
        RECT 76.760 -9.860 77.210 -9.770 ;
        RECT 79.610 -9.860 80.070 -9.780 ;
        RECT 76.760 -10.090 80.070 -9.860 ;
        RECT 76.760 -10.280 77.210 -10.090 ;
        RECT 79.610 -10.280 80.070 -10.090 ;
        RECT 76.760 -10.510 80.070 -10.280 ;
        RECT 76.760 -10.600 77.210 -10.510 ;
        RECT 79.610 -10.590 80.070 -10.510 ;
        RECT 83.560 -9.860 84.020 -9.780 ;
        RECT 86.420 -9.860 86.870 -9.770 ;
        RECT 83.560 -10.090 86.870 -9.860 ;
        RECT 83.560 -10.280 84.020 -10.090 ;
        RECT 86.420 -10.280 86.870 -10.090 ;
        RECT 83.560 -10.510 86.870 -10.280 ;
        RECT 83.560 -10.590 84.020 -10.510 ;
        RECT 86.420 -10.600 86.870 -10.510 ;
        RECT 90.260 -9.860 90.710 -9.770 ;
        RECT 93.110 -9.860 93.570 -9.780 ;
        RECT 90.260 -10.090 93.570 -9.860 ;
        RECT 90.260 -10.280 90.710 -10.090 ;
        RECT 93.110 -10.280 93.570 -10.090 ;
        RECT 90.260 -10.510 93.570 -10.280 ;
        RECT 90.260 -10.600 90.710 -10.510 ;
        RECT 93.110 -10.590 93.570 -10.510 ;
        RECT 97.060 -9.860 97.520 -9.780 ;
        RECT 99.920 -9.860 100.370 -9.770 ;
        RECT 97.060 -10.090 100.370 -9.860 ;
        RECT 97.060 -10.280 97.520 -10.090 ;
        RECT 99.920 -10.280 100.370 -10.090 ;
        RECT 97.060 -10.510 100.370 -10.280 ;
        RECT 97.060 -10.590 97.520 -10.510 ;
        RECT 99.920 -10.600 100.370 -10.510 ;
        RECT 103.760 -9.860 104.210 -9.770 ;
        RECT 106.610 -9.860 107.070 -9.780 ;
        RECT 103.760 -10.090 107.070 -9.860 ;
        RECT 103.760 -10.280 104.210 -10.090 ;
        RECT 106.610 -10.280 107.070 -10.090 ;
        RECT 103.760 -10.510 107.070 -10.280 ;
        RECT 103.760 -10.600 104.210 -10.510 ;
        RECT 106.610 -10.590 107.070 -10.510 ;
        RECT 110.560 -9.860 111.020 -9.780 ;
        RECT 113.420 -9.860 113.870 -9.770 ;
        RECT 110.560 -10.090 113.870 -9.860 ;
        RECT 110.560 -10.280 111.020 -10.090 ;
        RECT 113.420 -10.280 113.870 -10.090 ;
        RECT 110.560 -10.510 113.870 -10.280 ;
        RECT 110.560 -10.590 111.020 -10.510 ;
        RECT 113.420 -10.600 113.870 -10.510 ;
        RECT 117.260 -9.860 117.710 -9.770 ;
        RECT 120.110 -9.860 120.570 -9.780 ;
        RECT 117.260 -10.090 120.570 -9.860 ;
        RECT 117.260 -10.280 117.710 -10.090 ;
        RECT 120.110 -10.280 120.570 -10.090 ;
        RECT 117.260 -10.510 120.570 -10.280 ;
        RECT 117.260 -10.600 117.710 -10.510 ;
        RECT 120.110 -10.590 120.570 -10.510 ;
        RECT 124.060 -9.860 124.520 -9.780 ;
        RECT 126.920 -9.860 127.370 -9.770 ;
        RECT 124.060 -10.090 127.370 -9.860 ;
        RECT 124.060 -10.280 124.520 -10.090 ;
        RECT 126.920 -10.280 127.370 -10.090 ;
        RECT 124.060 -10.510 127.370 -10.280 ;
        RECT 124.060 -10.590 124.520 -10.510 ;
        RECT 126.920 -10.600 127.370 -10.510 ;
        RECT 130.760 -9.860 131.210 -9.770 ;
        RECT 133.610 -9.860 134.070 -9.780 ;
        RECT 130.760 -10.090 134.070 -9.860 ;
        RECT 130.760 -10.280 131.210 -10.090 ;
        RECT 133.610 -10.280 134.070 -10.090 ;
        RECT 130.760 -10.510 134.070 -10.280 ;
        RECT 130.760 -10.600 131.210 -10.510 ;
        RECT 133.610 -10.590 134.070 -10.510 ;
        RECT 137.560 -9.860 138.020 -9.780 ;
        RECT 140.420 -9.860 140.870 -9.770 ;
        RECT 137.560 -10.090 140.870 -9.860 ;
        RECT 137.560 -10.280 138.020 -10.090 ;
        RECT 140.420 -10.280 140.870 -10.090 ;
        RECT 137.560 -10.510 140.870 -10.280 ;
        RECT 137.560 -10.590 138.020 -10.510 ;
        RECT 140.420 -10.600 140.870 -10.510 ;
        RECT 144.260 -9.860 144.710 -9.770 ;
        RECT 147.110 -9.860 147.570 -9.780 ;
        RECT 144.260 -10.090 147.570 -9.860 ;
        RECT 144.260 -10.280 144.710 -10.090 ;
        RECT 147.110 -10.280 147.570 -10.090 ;
        RECT 144.260 -10.510 147.570 -10.280 ;
        RECT 144.260 -10.600 144.710 -10.510 ;
        RECT 147.110 -10.590 147.570 -10.510 ;
        RECT 151.060 -9.860 151.520 -9.780 ;
        RECT 153.920 -9.860 154.370 -9.770 ;
        RECT 151.060 -10.090 154.370 -9.860 ;
        RECT 151.060 -10.280 151.520 -10.090 ;
        RECT 153.920 -10.280 154.370 -10.090 ;
        RECT 151.060 -10.510 154.370 -10.280 ;
        RECT 151.060 -10.590 151.520 -10.510 ;
        RECT 153.920 -10.600 154.370 -10.510 ;
        RECT 157.760 -9.860 158.210 -9.770 ;
        RECT 160.610 -9.860 161.070 -9.780 ;
        RECT 157.760 -10.090 161.070 -9.860 ;
        RECT 157.760 -10.280 158.210 -10.090 ;
        RECT 160.610 -10.280 161.070 -10.090 ;
        RECT 157.760 -10.510 161.070 -10.280 ;
        RECT 157.760 -10.600 158.210 -10.510 ;
        RECT 160.610 -10.590 161.070 -10.510 ;
        RECT 164.560 -9.860 165.020 -9.780 ;
        RECT 167.420 -9.860 167.870 -9.770 ;
        RECT 164.560 -10.090 167.870 -9.860 ;
        RECT 164.560 -10.280 165.020 -10.090 ;
        RECT 167.420 -10.280 167.870 -10.090 ;
        RECT 164.560 -10.510 167.870 -10.280 ;
        RECT 164.560 -10.590 165.020 -10.510 ;
        RECT 167.420 -10.600 167.870 -10.510 ;
        RECT 171.260 -9.860 171.710 -9.770 ;
        RECT 174.110 -9.860 174.570 -9.780 ;
        RECT 171.260 -10.090 174.570 -9.860 ;
        RECT 171.260 -10.280 171.710 -10.090 ;
        RECT 174.110 -10.280 174.570 -10.090 ;
        RECT 171.260 -10.510 174.570 -10.280 ;
        RECT 171.260 -10.600 171.710 -10.510 ;
        RECT 174.110 -10.590 174.570 -10.510 ;
        RECT 178.060 -9.860 178.520 -9.780 ;
        RECT 180.920 -9.860 181.370 -9.770 ;
        RECT 178.060 -10.090 181.370 -9.860 ;
        RECT 178.060 -10.280 178.520 -10.090 ;
        RECT 180.920 -10.280 181.370 -10.090 ;
        RECT 178.060 -10.510 181.370 -10.280 ;
        RECT 178.060 -10.590 178.520 -10.510 ;
        RECT 180.920 -10.600 181.370 -10.510 ;
        RECT 184.760 -9.860 185.210 -9.770 ;
        RECT 187.610 -9.860 188.070 -9.780 ;
        RECT 184.760 -10.090 188.070 -9.860 ;
        RECT 184.760 -10.280 185.210 -10.090 ;
        RECT 187.610 -10.280 188.070 -10.090 ;
        RECT 184.760 -10.510 188.070 -10.280 ;
        RECT 184.760 -10.600 185.210 -10.510 ;
        RECT 187.610 -10.590 188.070 -10.510 ;
        RECT 191.560 -9.860 192.020 -9.780 ;
        RECT 194.420 -9.860 194.870 -9.770 ;
        RECT 191.560 -10.090 194.870 -9.860 ;
        RECT 191.560 -10.280 192.020 -10.090 ;
        RECT 194.420 -10.280 194.870 -10.090 ;
        RECT 191.560 -10.510 194.870 -10.280 ;
        RECT 191.560 -10.590 192.020 -10.510 ;
        RECT 194.420 -10.600 194.870 -10.510 ;
        RECT 198.260 -9.860 198.710 -9.770 ;
        RECT 201.110 -9.860 201.570 -9.780 ;
        RECT 198.260 -10.090 201.570 -9.860 ;
        RECT 198.260 -10.280 198.710 -10.090 ;
        RECT 201.110 -10.280 201.570 -10.090 ;
        RECT 198.260 -10.510 201.570 -10.280 ;
        RECT 198.260 -10.600 198.710 -10.510 ;
        RECT 201.110 -10.590 201.570 -10.510 ;
        RECT 205.060 -9.860 205.520 -9.780 ;
        RECT 207.920 -9.860 208.370 -9.770 ;
        RECT 205.060 -10.090 208.370 -9.860 ;
        RECT 205.060 -10.280 205.520 -10.090 ;
        RECT 207.920 -10.280 208.370 -10.090 ;
        RECT 205.060 -10.510 208.370 -10.280 ;
        RECT 205.060 -10.590 205.520 -10.510 ;
        RECT 207.920 -10.600 208.370 -10.510 ;
        RECT 211.760 -9.860 212.210 -9.770 ;
        RECT 214.610 -9.860 215.070 -9.780 ;
        RECT 211.760 -10.090 215.070 -9.860 ;
        RECT 211.760 -10.280 212.210 -10.090 ;
        RECT 214.610 -10.280 215.070 -10.090 ;
        RECT 211.760 -10.510 215.070 -10.280 ;
        RECT 211.760 -10.600 212.210 -10.510 ;
        RECT 214.610 -10.590 215.070 -10.510 ;
        RECT 9.260 -13.470 9.710 -13.380 ;
        RECT 12.110 -13.470 12.570 -13.390 ;
        RECT 9.260 -13.700 12.570 -13.470 ;
        RECT 9.260 -13.890 9.710 -13.700 ;
        RECT 12.110 -13.890 12.570 -13.700 ;
        RECT 9.260 -14.120 12.570 -13.890 ;
        RECT 9.260 -14.210 9.710 -14.120 ;
        RECT 12.110 -14.200 12.570 -14.120 ;
        RECT 16.060 -13.470 16.520 -13.390 ;
        RECT 18.920 -13.470 19.370 -13.380 ;
        RECT 16.060 -13.700 19.370 -13.470 ;
        RECT 16.060 -13.890 16.520 -13.700 ;
        RECT 18.920 -13.890 19.370 -13.700 ;
        RECT 16.060 -14.120 19.370 -13.890 ;
        RECT 16.060 -14.200 16.520 -14.120 ;
        RECT 18.920 -14.210 19.370 -14.120 ;
        RECT 22.760 -13.470 23.210 -13.380 ;
        RECT 25.610 -13.470 26.070 -13.390 ;
        RECT 22.760 -13.700 26.070 -13.470 ;
        RECT 22.760 -13.890 23.210 -13.700 ;
        RECT 25.610 -13.890 26.070 -13.700 ;
        RECT 22.760 -14.120 26.070 -13.890 ;
        RECT 22.760 -14.210 23.210 -14.120 ;
        RECT 25.610 -14.200 26.070 -14.120 ;
        RECT 29.560 -13.470 30.020 -13.390 ;
        RECT 32.420 -13.470 32.870 -13.380 ;
        RECT 29.560 -13.700 32.870 -13.470 ;
        RECT 29.560 -13.890 30.020 -13.700 ;
        RECT 32.420 -13.890 32.870 -13.700 ;
        RECT 29.560 -14.120 32.870 -13.890 ;
        RECT 29.560 -14.200 30.020 -14.120 ;
        RECT 32.420 -14.210 32.870 -14.120 ;
        RECT 36.260 -13.470 36.710 -13.380 ;
        RECT 39.110 -13.470 39.570 -13.390 ;
        RECT 36.260 -13.700 39.570 -13.470 ;
        RECT 36.260 -13.890 36.710 -13.700 ;
        RECT 39.110 -13.890 39.570 -13.700 ;
        RECT 36.260 -14.120 39.570 -13.890 ;
        RECT 36.260 -14.210 36.710 -14.120 ;
        RECT 39.110 -14.200 39.570 -14.120 ;
        RECT 43.060 -13.470 43.520 -13.390 ;
        RECT 45.920 -13.470 46.370 -13.380 ;
        RECT 43.060 -13.700 46.370 -13.470 ;
        RECT 43.060 -13.890 43.520 -13.700 ;
        RECT 45.920 -13.890 46.370 -13.700 ;
        RECT 43.060 -14.120 46.370 -13.890 ;
        RECT 43.060 -14.200 43.520 -14.120 ;
        RECT 45.920 -14.210 46.370 -14.120 ;
        RECT 49.760 -13.470 50.210 -13.380 ;
        RECT 52.610 -13.470 53.070 -13.390 ;
        RECT 49.760 -13.700 53.070 -13.470 ;
        RECT 49.760 -13.890 50.210 -13.700 ;
        RECT 52.610 -13.890 53.070 -13.700 ;
        RECT 49.760 -14.120 53.070 -13.890 ;
        RECT 49.760 -14.210 50.210 -14.120 ;
        RECT 52.610 -14.200 53.070 -14.120 ;
        RECT 56.560 -13.470 57.020 -13.390 ;
        RECT 59.420 -13.470 59.870 -13.380 ;
        RECT 56.560 -13.700 59.870 -13.470 ;
        RECT 56.560 -13.890 57.020 -13.700 ;
        RECT 59.420 -13.890 59.870 -13.700 ;
        RECT 56.560 -14.120 59.870 -13.890 ;
        RECT 56.560 -14.200 57.020 -14.120 ;
        RECT 59.420 -14.210 59.870 -14.120 ;
        RECT 63.260 -13.470 63.710 -13.380 ;
        RECT 66.110 -13.470 66.570 -13.390 ;
        RECT 63.260 -13.700 66.570 -13.470 ;
        RECT 63.260 -13.890 63.710 -13.700 ;
        RECT 66.110 -13.890 66.570 -13.700 ;
        RECT 63.260 -14.120 66.570 -13.890 ;
        RECT 63.260 -14.210 63.710 -14.120 ;
        RECT 66.110 -14.200 66.570 -14.120 ;
        RECT 70.060 -13.470 70.520 -13.390 ;
        RECT 72.920 -13.470 73.370 -13.380 ;
        RECT 70.060 -13.700 73.370 -13.470 ;
        RECT 70.060 -13.890 70.520 -13.700 ;
        RECT 72.920 -13.890 73.370 -13.700 ;
        RECT 70.060 -14.120 73.370 -13.890 ;
        RECT 70.060 -14.200 70.520 -14.120 ;
        RECT 72.920 -14.210 73.370 -14.120 ;
        RECT 76.760 -13.470 77.210 -13.380 ;
        RECT 79.610 -13.470 80.070 -13.390 ;
        RECT 76.760 -13.700 80.070 -13.470 ;
        RECT 76.760 -13.890 77.210 -13.700 ;
        RECT 79.610 -13.890 80.070 -13.700 ;
        RECT 76.760 -14.120 80.070 -13.890 ;
        RECT 76.760 -14.210 77.210 -14.120 ;
        RECT 79.610 -14.200 80.070 -14.120 ;
        RECT 83.560 -13.470 84.020 -13.390 ;
        RECT 86.420 -13.470 86.870 -13.380 ;
        RECT 83.560 -13.700 86.870 -13.470 ;
        RECT 83.560 -13.890 84.020 -13.700 ;
        RECT 86.420 -13.890 86.870 -13.700 ;
        RECT 83.560 -14.120 86.870 -13.890 ;
        RECT 83.560 -14.200 84.020 -14.120 ;
        RECT 86.420 -14.210 86.870 -14.120 ;
        RECT 90.260 -13.470 90.710 -13.380 ;
        RECT 93.110 -13.470 93.570 -13.390 ;
        RECT 90.260 -13.700 93.570 -13.470 ;
        RECT 90.260 -13.890 90.710 -13.700 ;
        RECT 93.110 -13.890 93.570 -13.700 ;
        RECT 90.260 -14.120 93.570 -13.890 ;
        RECT 90.260 -14.210 90.710 -14.120 ;
        RECT 93.110 -14.200 93.570 -14.120 ;
        RECT 97.060 -13.470 97.520 -13.390 ;
        RECT 99.920 -13.470 100.370 -13.380 ;
        RECT 97.060 -13.700 100.370 -13.470 ;
        RECT 97.060 -13.890 97.520 -13.700 ;
        RECT 99.920 -13.890 100.370 -13.700 ;
        RECT 97.060 -14.120 100.370 -13.890 ;
        RECT 97.060 -14.200 97.520 -14.120 ;
        RECT 99.920 -14.210 100.370 -14.120 ;
        RECT 103.760 -13.470 104.210 -13.380 ;
        RECT 106.610 -13.470 107.070 -13.390 ;
        RECT 103.760 -13.700 107.070 -13.470 ;
        RECT 103.760 -13.890 104.210 -13.700 ;
        RECT 106.610 -13.890 107.070 -13.700 ;
        RECT 103.760 -14.120 107.070 -13.890 ;
        RECT 103.760 -14.210 104.210 -14.120 ;
        RECT 106.610 -14.200 107.070 -14.120 ;
        RECT 110.560 -13.470 111.020 -13.390 ;
        RECT 113.420 -13.470 113.870 -13.380 ;
        RECT 110.560 -13.700 113.870 -13.470 ;
        RECT 110.560 -13.890 111.020 -13.700 ;
        RECT 113.420 -13.890 113.870 -13.700 ;
        RECT 110.560 -14.120 113.870 -13.890 ;
        RECT 110.560 -14.200 111.020 -14.120 ;
        RECT 113.420 -14.210 113.870 -14.120 ;
        RECT 117.260 -13.470 117.710 -13.380 ;
        RECT 120.110 -13.470 120.570 -13.390 ;
        RECT 117.260 -13.700 120.570 -13.470 ;
        RECT 117.260 -13.890 117.710 -13.700 ;
        RECT 120.110 -13.890 120.570 -13.700 ;
        RECT 117.260 -14.120 120.570 -13.890 ;
        RECT 117.260 -14.210 117.710 -14.120 ;
        RECT 120.110 -14.200 120.570 -14.120 ;
        RECT 124.060 -13.470 124.520 -13.390 ;
        RECT 126.920 -13.470 127.370 -13.380 ;
        RECT 124.060 -13.700 127.370 -13.470 ;
        RECT 124.060 -13.890 124.520 -13.700 ;
        RECT 126.920 -13.890 127.370 -13.700 ;
        RECT 124.060 -14.120 127.370 -13.890 ;
        RECT 124.060 -14.200 124.520 -14.120 ;
        RECT 126.920 -14.210 127.370 -14.120 ;
        RECT 130.760 -13.470 131.210 -13.380 ;
        RECT 133.610 -13.470 134.070 -13.390 ;
        RECT 130.760 -13.700 134.070 -13.470 ;
        RECT 130.760 -13.890 131.210 -13.700 ;
        RECT 133.610 -13.890 134.070 -13.700 ;
        RECT 130.760 -14.120 134.070 -13.890 ;
        RECT 130.760 -14.210 131.210 -14.120 ;
        RECT 133.610 -14.200 134.070 -14.120 ;
        RECT 137.560 -13.470 138.020 -13.390 ;
        RECT 140.420 -13.470 140.870 -13.380 ;
        RECT 137.560 -13.700 140.870 -13.470 ;
        RECT 137.560 -13.890 138.020 -13.700 ;
        RECT 140.420 -13.890 140.870 -13.700 ;
        RECT 137.560 -14.120 140.870 -13.890 ;
        RECT 137.560 -14.200 138.020 -14.120 ;
        RECT 140.420 -14.210 140.870 -14.120 ;
        RECT 144.260 -13.470 144.710 -13.380 ;
        RECT 147.110 -13.470 147.570 -13.390 ;
        RECT 144.260 -13.700 147.570 -13.470 ;
        RECT 144.260 -13.890 144.710 -13.700 ;
        RECT 147.110 -13.890 147.570 -13.700 ;
        RECT 144.260 -14.120 147.570 -13.890 ;
        RECT 144.260 -14.210 144.710 -14.120 ;
        RECT 147.110 -14.200 147.570 -14.120 ;
        RECT 151.060 -13.470 151.520 -13.390 ;
        RECT 153.920 -13.470 154.370 -13.380 ;
        RECT 151.060 -13.700 154.370 -13.470 ;
        RECT 151.060 -13.890 151.520 -13.700 ;
        RECT 153.920 -13.890 154.370 -13.700 ;
        RECT 151.060 -14.120 154.370 -13.890 ;
        RECT 151.060 -14.200 151.520 -14.120 ;
        RECT 153.920 -14.210 154.370 -14.120 ;
        RECT 157.760 -13.470 158.210 -13.380 ;
        RECT 160.610 -13.470 161.070 -13.390 ;
        RECT 157.760 -13.700 161.070 -13.470 ;
        RECT 157.760 -13.890 158.210 -13.700 ;
        RECT 160.610 -13.890 161.070 -13.700 ;
        RECT 157.760 -14.120 161.070 -13.890 ;
        RECT 157.760 -14.210 158.210 -14.120 ;
        RECT 160.610 -14.200 161.070 -14.120 ;
        RECT 164.560 -13.470 165.020 -13.390 ;
        RECT 167.420 -13.470 167.870 -13.380 ;
        RECT 164.560 -13.700 167.870 -13.470 ;
        RECT 164.560 -13.890 165.020 -13.700 ;
        RECT 167.420 -13.890 167.870 -13.700 ;
        RECT 164.560 -14.120 167.870 -13.890 ;
        RECT 164.560 -14.200 165.020 -14.120 ;
        RECT 167.420 -14.210 167.870 -14.120 ;
        RECT 171.260 -13.470 171.710 -13.380 ;
        RECT 174.110 -13.470 174.570 -13.390 ;
        RECT 171.260 -13.700 174.570 -13.470 ;
        RECT 171.260 -13.890 171.710 -13.700 ;
        RECT 174.110 -13.890 174.570 -13.700 ;
        RECT 171.260 -14.120 174.570 -13.890 ;
        RECT 171.260 -14.210 171.710 -14.120 ;
        RECT 174.110 -14.200 174.570 -14.120 ;
        RECT 178.060 -13.470 178.520 -13.390 ;
        RECT 180.920 -13.470 181.370 -13.380 ;
        RECT 178.060 -13.700 181.370 -13.470 ;
        RECT 178.060 -13.890 178.520 -13.700 ;
        RECT 180.920 -13.890 181.370 -13.700 ;
        RECT 178.060 -14.120 181.370 -13.890 ;
        RECT 178.060 -14.200 178.520 -14.120 ;
        RECT 180.920 -14.210 181.370 -14.120 ;
        RECT 184.760 -13.470 185.210 -13.380 ;
        RECT 187.610 -13.470 188.070 -13.390 ;
        RECT 184.760 -13.700 188.070 -13.470 ;
        RECT 184.760 -13.890 185.210 -13.700 ;
        RECT 187.610 -13.890 188.070 -13.700 ;
        RECT 184.760 -14.120 188.070 -13.890 ;
        RECT 184.760 -14.210 185.210 -14.120 ;
        RECT 187.610 -14.200 188.070 -14.120 ;
        RECT 191.560 -13.470 192.020 -13.390 ;
        RECT 194.420 -13.470 194.870 -13.380 ;
        RECT 191.560 -13.700 194.870 -13.470 ;
        RECT 191.560 -13.890 192.020 -13.700 ;
        RECT 194.420 -13.890 194.870 -13.700 ;
        RECT 191.560 -14.120 194.870 -13.890 ;
        RECT 191.560 -14.200 192.020 -14.120 ;
        RECT 194.420 -14.210 194.870 -14.120 ;
        RECT 198.260 -13.470 198.710 -13.380 ;
        RECT 201.110 -13.470 201.570 -13.390 ;
        RECT 198.260 -13.700 201.570 -13.470 ;
        RECT 198.260 -13.890 198.710 -13.700 ;
        RECT 201.110 -13.890 201.570 -13.700 ;
        RECT 198.260 -14.120 201.570 -13.890 ;
        RECT 198.260 -14.210 198.710 -14.120 ;
        RECT 201.110 -14.200 201.570 -14.120 ;
        RECT 205.060 -13.470 205.520 -13.390 ;
        RECT 207.920 -13.470 208.370 -13.380 ;
        RECT 205.060 -13.700 208.370 -13.470 ;
        RECT 205.060 -13.890 205.520 -13.700 ;
        RECT 207.920 -13.890 208.370 -13.700 ;
        RECT 205.060 -14.120 208.370 -13.890 ;
        RECT 205.060 -14.200 205.520 -14.120 ;
        RECT 207.920 -14.210 208.370 -14.120 ;
        RECT 211.760 -13.470 212.210 -13.380 ;
        RECT 214.610 -13.470 215.070 -13.390 ;
        RECT 211.760 -13.700 215.070 -13.470 ;
        RECT 211.760 -13.890 212.210 -13.700 ;
        RECT 214.610 -13.890 215.070 -13.700 ;
        RECT 211.760 -14.120 215.070 -13.890 ;
        RECT 211.760 -14.210 212.210 -14.120 ;
        RECT 214.610 -14.200 215.070 -14.120 ;
        RECT 9.260 -17.080 9.710 -16.990 ;
        RECT 12.110 -17.080 12.570 -17.000 ;
        RECT 9.260 -17.310 12.570 -17.080 ;
        RECT 9.260 -17.500 9.710 -17.310 ;
        RECT 12.110 -17.500 12.570 -17.310 ;
        RECT 9.260 -17.730 12.570 -17.500 ;
        RECT 9.260 -17.820 9.710 -17.730 ;
        RECT 12.110 -17.810 12.570 -17.730 ;
        RECT 16.060 -17.080 16.520 -17.000 ;
        RECT 18.920 -17.080 19.370 -16.990 ;
        RECT 16.060 -17.310 19.370 -17.080 ;
        RECT 16.060 -17.500 16.520 -17.310 ;
        RECT 18.920 -17.500 19.370 -17.310 ;
        RECT 16.060 -17.730 19.370 -17.500 ;
        RECT 16.060 -17.810 16.520 -17.730 ;
        RECT 18.920 -17.820 19.370 -17.730 ;
        RECT 22.760 -17.080 23.210 -16.990 ;
        RECT 25.610 -17.080 26.070 -17.000 ;
        RECT 22.760 -17.310 26.070 -17.080 ;
        RECT 22.760 -17.500 23.210 -17.310 ;
        RECT 25.610 -17.500 26.070 -17.310 ;
        RECT 22.760 -17.730 26.070 -17.500 ;
        RECT 22.760 -17.820 23.210 -17.730 ;
        RECT 25.610 -17.810 26.070 -17.730 ;
        RECT 29.560 -17.080 30.020 -17.000 ;
        RECT 32.420 -17.080 32.870 -16.990 ;
        RECT 29.560 -17.310 32.870 -17.080 ;
        RECT 29.560 -17.500 30.020 -17.310 ;
        RECT 32.420 -17.500 32.870 -17.310 ;
        RECT 29.560 -17.730 32.870 -17.500 ;
        RECT 29.560 -17.810 30.020 -17.730 ;
        RECT 32.420 -17.820 32.870 -17.730 ;
        RECT 36.260 -17.080 36.710 -16.990 ;
        RECT 39.110 -17.080 39.570 -17.000 ;
        RECT 36.260 -17.310 39.570 -17.080 ;
        RECT 36.260 -17.500 36.710 -17.310 ;
        RECT 39.110 -17.500 39.570 -17.310 ;
        RECT 36.260 -17.730 39.570 -17.500 ;
        RECT 36.260 -17.820 36.710 -17.730 ;
        RECT 39.110 -17.810 39.570 -17.730 ;
        RECT 43.060 -17.080 43.520 -17.000 ;
        RECT 45.920 -17.080 46.370 -16.990 ;
        RECT 43.060 -17.310 46.370 -17.080 ;
        RECT 43.060 -17.500 43.520 -17.310 ;
        RECT 45.920 -17.500 46.370 -17.310 ;
        RECT 43.060 -17.730 46.370 -17.500 ;
        RECT 43.060 -17.810 43.520 -17.730 ;
        RECT 45.920 -17.820 46.370 -17.730 ;
        RECT 49.760 -17.080 50.210 -16.990 ;
        RECT 52.610 -17.080 53.070 -17.000 ;
        RECT 49.760 -17.310 53.070 -17.080 ;
        RECT 49.760 -17.500 50.210 -17.310 ;
        RECT 52.610 -17.500 53.070 -17.310 ;
        RECT 49.760 -17.730 53.070 -17.500 ;
        RECT 49.760 -17.820 50.210 -17.730 ;
        RECT 52.610 -17.810 53.070 -17.730 ;
        RECT 56.560 -17.080 57.020 -17.000 ;
        RECT 59.420 -17.080 59.870 -16.990 ;
        RECT 56.560 -17.310 59.870 -17.080 ;
        RECT 56.560 -17.500 57.020 -17.310 ;
        RECT 59.420 -17.500 59.870 -17.310 ;
        RECT 56.560 -17.730 59.870 -17.500 ;
        RECT 56.560 -17.810 57.020 -17.730 ;
        RECT 59.420 -17.820 59.870 -17.730 ;
        RECT 63.260 -17.080 63.710 -16.990 ;
        RECT 66.110 -17.080 66.570 -17.000 ;
        RECT 63.260 -17.310 66.570 -17.080 ;
        RECT 63.260 -17.500 63.710 -17.310 ;
        RECT 66.110 -17.500 66.570 -17.310 ;
        RECT 63.260 -17.730 66.570 -17.500 ;
        RECT 63.260 -17.820 63.710 -17.730 ;
        RECT 66.110 -17.810 66.570 -17.730 ;
        RECT 70.060 -17.080 70.520 -17.000 ;
        RECT 72.920 -17.080 73.370 -16.990 ;
        RECT 70.060 -17.310 73.370 -17.080 ;
        RECT 70.060 -17.500 70.520 -17.310 ;
        RECT 72.920 -17.500 73.370 -17.310 ;
        RECT 70.060 -17.730 73.370 -17.500 ;
        RECT 70.060 -17.810 70.520 -17.730 ;
        RECT 72.920 -17.820 73.370 -17.730 ;
        RECT 76.760 -17.080 77.210 -16.990 ;
        RECT 79.610 -17.080 80.070 -17.000 ;
        RECT 76.760 -17.310 80.070 -17.080 ;
        RECT 76.760 -17.500 77.210 -17.310 ;
        RECT 79.610 -17.500 80.070 -17.310 ;
        RECT 76.760 -17.730 80.070 -17.500 ;
        RECT 76.760 -17.820 77.210 -17.730 ;
        RECT 79.610 -17.810 80.070 -17.730 ;
        RECT 83.560 -17.080 84.020 -17.000 ;
        RECT 86.420 -17.080 86.870 -16.990 ;
        RECT 83.560 -17.310 86.870 -17.080 ;
        RECT 83.560 -17.500 84.020 -17.310 ;
        RECT 86.420 -17.500 86.870 -17.310 ;
        RECT 83.560 -17.730 86.870 -17.500 ;
        RECT 83.560 -17.810 84.020 -17.730 ;
        RECT 86.420 -17.820 86.870 -17.730 ;
        RECT 90.260 -17.080 90.710 -16.990 ;
        RECT 93.110 -17.080 93.570 -17.000 ;
        RECT 90.260 -17.310 93.570 -17.080 ;
        RECT 90.260 -17.500 90.710 -17.310 ;
        RECT 93.110 -17.500 93.570 -17.310 ;
        RECT 90.260 -17.730 93.570 -17.500 ;
        RECT 90.260 -17.820 90.710 -17.730 ;
        RECT 93.110 -17.810 93.570 -17.730 ;
        RECT 97.060 -17.080 97.520 -17.000 ;
        RECT 99.920 -17.080 100.370 -16.990 ;
        RECT 97.060 -17.310 100.370 -17.080 ;
        RECT 97.060 -17.500 97.520 -17.310 ;
        RECT 99.920 -17.500 100.370 -17.310 ;
        RECT 97.060 -17.730 100.370 -17.500 ;
        RECT 97.060 -17.810 97.520 -17.730 ;
        RECT 99.920 -17.820 100.370 -17.730 ;
        RECT 103.760 -17.080 104.210 -16.990 ;
        RECT 106.610 -17.080 107.070 -17.000 ;
        RECT 103.760 -17.310 107.070 -17.080 ;
        RECT 103.760 -17.500 104.210 -17.310 ;
        RECT 106.610 -17.500 107.070 -17.310 ;
        RECT 103.760 -17.730 107.070 -17.500 ;
        RECT 103.760 -17.820 104.210 -17.730 ;
        RECT 106.610 -17.810 107.070 -17.730 ;
        RECT 110.560 -17.080 111.020 -17.000 ;
        RECT 113.420 -17.080 113.870 -16.990 ;
        RECT 110.560 -17.310 113.870 -17.080 ;
        RECT 110.560 -17.500 111.020 -17.310 ;
        RECT 113.420 -17.500 113.870 -17.310 ;
        RECT 110.560 -17.730 113.870 -17.500 ;
        RECT 110.560 -17.810 111.020 -17.730 ;
        RECT 113.420 -17.820 113.870 -17.730 ;
        RECT 117.260 -17.080 117.710 -16.990 ;
        RECT 120.110 -17.080 120.570 -17.000 ;
        RECT 117.260 -17.310 120.570 -17.080 ;
        RECT 117.260 -17.500 117.710 -17.310 ;
        RECT 120.110 -17.500 120.570 -17.310 ;
        RECT 117.260 -17.730 120.570 -17.500 ;
        RECT 117.260 -17.820 117.710 -17.730 ;
        RECT 120.110 -17.810 120.570 -17.730 ;
        RECT 124.060 -17.080 124.520 -17.000 ;
        RECT 126.920 -17.080 127.370 -16.990 ;
        RECT 124.060 -17.310 127.370 -17.080 ;
        RECT 124.060 -17.500 124.520 -17.310 ;
        RECT 126.920 -17.500 127.370 -17.310 ;
        RECT 124.060 -17.730 127.370 -17.500 ;
        RECT 124.060 -17.810 124.520 -17.730 ;
        RECT 126.920 -17.820 127.370 -17.730 ;
        RECT 130.760 -17.080 131.210 -16.990 ;
        RECT 133.610 -17.080 134.070 -17.000 ;
        RECT 130.760 -17.310 134.070 -17.080 ;
        RECT 130.760 -17.500 131.210 -17.310 ;
        RECT 133.610 -17.500 134.070 -17.310 ;
        RECT 130.760 -17.730 134.070 -17.500 ;
        RECT 130.760 -17.820 131.210 -17.730 ;
        RECT 133.610 -17.810 134.070 -17.730 ;
        RECT 137.560 -17.080 138.020 -17.000 ;
        RECT 140.420 -17.080 140.870 -16.990 ;
        RECT 137.560 -17.310 140.870 -17.080 ;
        RECT 137.560 -17.500 138.020 -17.310 ;
        RECT 140.420 -17.500 140.870 -17.310 ;
        RECT 137.560 -17.730 140.870 -17.500 ;
        RECT 137.560 -17.810 138.020 -17.730 ;
        RECT 140.420 -17.820 140.870 -17.730 ;
        RECT 144.260 -17.080 144.710 -16.990 ;
        RECT 147.110 -17.080 147.570 -17.000 ;
        RECT 144.260 -17.310 147.570 -17.080 ;
        RECT 144.260 -17.500 144.710 -17.310 ;
        RECT 147.110 -17.500 147.570 -17.310 ;
        RECT 144.260 -17.730 147.570 -17.500 ;
        RECT 144.260 -17.820 144.710 -17.730 ;
        RECT 147.110 -17.810 147.570 -17.730 ;
        RECT 151.060 -17.080 151.520 -17.000 ;
        RECT 153.920 -17.080 154.370 -16.990 ;
        RECT 151.060 -17.310 154.370 -17.080 ;
        RECT 151.060 -17.500 151.520 -17.310 ;
        RECT 153.920 -17.500 154.370 -17.310 ;
        RECT 151.060 -17.730 154.370 -17.500 ;
        RECT 151.060 -17.810 151.520 -17.730 ;
        RECT 153.920 -17.820 154.370 -17.730 ;
        RECT 157.760 -17.080 158.210 -16.990 ;
        RECT 160.610 -17.080 161.070 -17.000 ;
        RECT 157.760 -17.310 161.070 -17.080 ;
        RECT 157.760 -17.500 158.210 -17.310 ;
        RECT 160.610 -17.500 161.070 -17.310 ;
        RECT 157.760 -17.730 161.070 -17.500 ;
        RECT 157.760 -17.820 158.210 -17.730 ;
        RECT 160.610 -17.810 161.070 -17.730 ;
        RECT 164.560 -17.080 165.020 -17.000 ;
        RECT 167.420 -17.080 167.870 -16.990 ;
        RECT 164.560 -17.310 167.870 -17.080 ;
        RECT 164.560 -17.500 165.020 -17.310 ;
        RECT 167.420 -17.500 167.870 -17.310 ;
        RECT 164.560 -17.730 167.870 -17.500 ;
        RECT 164.560 -17.810 165.020 -17.730 ;
        RECT 167.420 -17.820 167.870 -17.730 ;
        RECT 171.260 -17.080 171.710 -16.990 ;
        RECT 174.110 -17.080 174.570 -17.000 ;
        RECT 171.260 -17.310 174.570 -17.080 ;
        RECT 171.260 -17.500 171.710 -17.310 ;
        RECT 174.110 -17.500 174.570 -17.310 ;
        RECT 171.260 -17.730 174.570 -17.500 ;
        RECT 171.260 -17.820 171.710 -17.730 ;
        RECT 174.110 -17.810 174.570 -17.730 ;
        RECT 178.060 -17.080 178.520 -17.000 ;
        RECT 180.920 -17.080 181.370 -16.990 ;
        RECT 178.060 -17.310 181.370 -17.080 ;
        RECT 178.060 -17.500 178.520 -17.310 ;
        RECT 180.920 -17.500 181.370 -17.310 ;
        RECT 178.060 -17.730 181.370 -17.500 ;
        RECT 178.060 -17.810 178.520 -17.730 ;
        RECT 180.920 -17.820 181.370 -17.730 ;
        RECT 184.760 -17.080 185.210 -16.990 ;
        RECT 187.610 -17.080 188.070 -17.000 ;
        RECT 184.760 -17.310 188.070 -17.080 ;
        RECT 184.760 -17.500 185.210 -17.310 ;
        RECT 187.610 -17.500 188.070 -17.310 ;
        RECT 184.760 -17.730 188.070 -17.500 ;
        RECT 184.760 -17.820 185.210 -17.730 ;
        RECT 187.610 -17.810 188.070 -17.730 ;
        RECT 191.560 -17.080 192.020 -17.000 ;
        RECT 194.420 -17.080 194.870 -16.990 ;
        RECT 191.560 -17.310 194.870 -17.080 ;
        RECT 191.560 -17.500 192.020 -17.310 ;
        RECT 194.420 -17.500 194.870 -17.310 ;
        RECT 191.560 -17.730 194.870 -17.500 ;
        RECT 191.560 -17.810 192.020 -17.730 ;
        RECT 194.420 -17.820 194.870 -17.730 ;
        RECT 198.260 -17.080 198.710 -16.990 ;
        RECT 201.110 -17.080 201.570 -17.000 ;
        RECT 198.260 -17.310 201.570 -17.080 ;
        RECT 198.260 -17.500 198.710 -17.310 ;
        RECT 201.110 -17.500 201.570 -17.310 ;
        RECT 198.260 -17.730 201.570 -17.500 ;
        RECT 198.260 -17.820 198.710 -17.730 ;
        RECT 201.110 -17.810 201.570 -17.730 ;
        RECT 205.060 -17.080 205.520 -17.000 ;
        RECT 207.920 -17.080 208.370 -16.990 ;
        RECT 205.060 -17.310 208.370 -17.080 ;
        RECT 205.060 -17.500 205.520 -17.310 ;
        RECT 207.920 -17.500 208.370 -17.310 ;
        RECT 205.060 -17.730 208.370 -17.500 ;
        RECT 205.060 -17.810 205.520 -17.730 ;
        RECT 207.920 -17.820 208.370 -17.730 ;
        RECT 211.760 -17.080 212.210 -16.990 ;
        RECT 214.610 -17.080 215.070 -17.000 ;
        RECT 211.760 -17.310 215.070 -17.080 ;
        RECT 211.760 -17.500 212.210 -17.310 ;
        RECT 214.610 -17.500 215.070 -17.310 ;
        RECT 211.760 -17.730 215.070 -17.500 ;
        RECT 211.760 -17.820 212.210 -17.730 ;
        RECT 214.610 -17.810 215.070 -17.730 ;
        RECT 9.260 -20.690 9.710 -20.600 ;
        RECT 12.110 -20.690 12.570 -20.610 ;
        RECT 9.260 -20.920 12.570 -20.690 ;
        RECT 9.260 -21.110 9.710 -20.920 ;
        RECT 12.110 -21.110 12.570 -20.920 ;
        RECT 9.260 -21.340 12.570 -21.110 ;
        RECT 9.260 -21.430 9.710 -21.340 ;
        RECT 12.110 -21.420 12.570 -21.340 ;
        RECT 16.060 -20.690 16.520 -20.610 ;
        RECT 18.920 -20.690 19.370 -20.600 ;
        RECT 16.060 -20.920 19.370 -20.690 ;
        RECT 16.060 -21.110 16.520 -20.920 ;
        RECT 18.920 -21.110 19.370 -20.920 ;
        RECT 16.060 -21.340 19.370 -21.110 ;
        RECT 16.060 -21.420 16.520 -21.340 ;
        RECT 18.920 -21.430 19.370 -21.340 ;
        RECT 22.760 -20.690 23.210 -20.600 ;
        RECT 25.610 -20.690 26.070 -20.610 ;
        RECT 22.760 -20.920 26.070 -20.690 ;
        RECT 22.760 -21.110 23.210 -20.920 ;
        RECT 25.610 -21.110 26.070 -20.920 ;
        RECT 22.760 -21.340 26.070 -21.110 ;
        RECT 22.760 -21.430 23.210 -21.340 ;
        RECT 25.610 -21.420 26.070 -21.340 ;
        RECT 29.560 -20.690 30.020 -20.610 ;
        RECT 32.420 -20.690 32.870 -20.600 ;
        RECT 29.560 -20.920 32.870 -20.690 ;
        RECT 29.560 -21.110 30.020 -20.920 ;
        RECT 32.420 -21.110 32.870 -20.920 ;
        RECT 29.560 -21.340 32.870 -21.110 ;
        RECT 29.560 -21.420 30.020 -21.340 ;
        RECT 32.420 -21.430 32.870 -21.340 ;
        RECT 36.260 -20.690 36.710 -20.600 ;
        RECT 39.110 -20.690 39.570 -20.610 ;
        RECT 36.260 -20.920 39.570 -20.690 ;
        RECT 36.260 -21.110 36.710 -20.920 ;
        RECT 39.110 -21.110 39.570 -20.920 ;
        RECT 36.260 -21.340 39.570 -21.110 ;
        RECT 36.260 -21.430 36.710 -21.340 ;
        RECT 39.110 -21.420 39.570 -21.340 ;
        RECT 43.060 -20.690 43.520 -20.610 ;
        RECT 45.920 -20.690 46.370 -20.600 ;
        RECT 43.060 -20.920 46.370 -20.690 ;
        RECT 43.060 -21.110 43.520 -20.920 ;
        RECT 45.920 -21.110 46.370 -20.920 ;
        RECT 43.060 -21.340 46.370 -21.110 ;
        RECT 43.060 -21.420 43.520 -21.340 ;
        RECT 45.920 -21.430 46.370 -21.340 ;
        RECT 49.760 -20.690 50.210 -20.600 ;
        RECT 52.610 -20.690 53.070 -20.610 ;
        RECT 49.760 -20.920 53.070 -20.690 ;
        RECT 49.760 -21.110 50.210 -20.920 ;
        RECT 52.610 -21.110 53.070 -20.920 ;
        RECT 49.760 -21.340 53.070 -21.110 ;
        RECT 49.760 -21.430 50.210 -21.340 ;
        RECT 52.610 -21.420 53.070 -21.340 ;
        RECT 56.560 -20.690 57.020 -20.610 ;
        RECT 59.420 -20.690 59.870 -20.600 ;
        RECT 56.560 -20.920 59.870 -20.690 ;
        RECT 56.560 -21.110 57.020 -20.920 ;
        RECT 59.420 -21.110 59.870 -20.920 ;
        RECT 56.560 -21.340 59.870 -21.110 ;
        RECT 56.560 -21.420 57.020 -21.340 ;
        RECT 59.420 -21.430 59.870 -21.340 ;
        RECT 63.260 -20.690 63.710 -20.600 ;
        RECT 66.110 -20.690 66.570 -20.610 ;
        RECT 63.260 -20.920 66.570 -20.690 ;
        RECT 63.260 -21.110 63.710 -20.920 ;
        RECT 66.110 -21.110 66.570 -20.920 ;
        RECT 63.260 -21.340 66.570 -21.110 ;
        RECT 63.260 -21.430 63.710 -21.340 ;
        RECT 66.110 -21.420 66.570 -21.340 ;
        RECT 70.060 -20.690 70.520 -20.610 ;
        RECT 72.920 -20.690 73.370 -20.600 ;
        RECT 70.060 -20.920 73.370 -20.690 ;
        RECT 70.060 -21.110 70.520 -20.920 ;
        RECT 72.920 -21.110 73.370 -20.920 ;
        RECT 70.060 -21.340 73.370 -21.110 ;
        RECT 70.060 -21.420 70.520 -21.340 ;
        RECT 72.920 -21.430 73.370 -21.340 ;
        RECT 76.760 -20.690 77.210 -20.600 ;
        RECT 79.610 -20.690 80.070 -20.610 ;
        RECT 76.760 -20.920 80.070 -20.690 ;
        RECT 76.760 -21.110 77.210 -20.920 ;
        RECT 79.610 -21.110 80.070 -20.920 ;
        RECT 76.760 -21.340 80.070 -21.110 ;
        RECT 76.760 -21.430 77.210 -21.340 ;
        RECT 79.610 -21.420 80.070 -21.340 ;
        RECT 83.560 -20.690 84.020 -20.610 ;
        RECT 86.420 -20.690 86.870 -20.600 ;
        RECT 83.560 -20.920 86.870 -20.690 ;
        RECT 83.560 -21.110 84.020 -20.920 ;
        RECT 86.420 -21.110 86.870 -20.920 ;
        RECT 83.560 -21.340 86.870 -21.110 ;
        RECT 83.560 -21.420 84.020 -21.340 ;
        RECT 86.420 -21.430 86.870 -21.340 ;
        RECT 90.260 -20.690 90.710 -20.600 ;
        RECT 93.110 -20.690 93.570 -20.610 ;
        RECT 90.260 -20.920 93.570 -20.690 ;
        RECT 90.260 -21.110 90.710 -20.920 ;
        RECT 93.110 -21.110 93.570 -20.920 ;
        RECT 90.260 -21.340 93.570 -21.110 ;
        RECT 90.260 -21.430 90.710 -21.340 ;
        RECT 93.110 -21.420 93.570 -21.340 ;
        RECT 97.060 -20.690 97.520 -20.610 ;
        RECT 99.920 -20.690 100.370 -20.600 ;
        RECT 97.060 -20.920 100.370 -20.690 ;
        RECT 97.060 -21.110 97.520 -20.920 ;
        RECT 99.920 -21.110 100.370 -20.920 ;
        RECT 97.060 -21.340 100.370 -21.110 ;
        RECT 97.060 -21.420 97.520 -21.340 ;
        RECT 99.920 -21.430 100.370 -21.340 ;
        RECT 103.760 -20.690 104.210 -20.600 ;
        RECT 106.610 -20.690 107.070 -20.610 ;
        RECT 103.760 -20.920 107.070 -20.690 ;
        RECT 103.760 -21.110 104.210 -20.920 ;
        RECT 106.610 -21.110 107.070 -20.920 ;
        RECT 103.760 -21.340 107.070 -21.110 ;
        RECT 103.760 -21.430 104.210 -21.340 ;
        RECT 106.610 -21.420 107.070 -21.340 ;
        RECT 110.560 -20.690 111.020 -20.610 ;
        RECT 113.420 -20.690 113.870 -20.600 ;
        RECT 110.560 -20.920 113.870 -20.690 ;
        RECT 110.560 -21.110 111.020 -20.920 ;
        RECT 113.420 -21.110 113.870 -20.920 ;
        RECT 110.560 -21.340 113.870 -21.110 ;
        RECT 110.560 -21.420 111.020 -21.340 ;
        RECT 113.420 -21.430 113.870 -21.340 ;
        RECT 117.260 -20.690 117.710 -20.600 ;
        RECT 120.110 -20.690 120.570 -20.610 ;
        RECT 117.260 -20.920 120.570 -20.690 ;
        RECT 117.260 -21.110 117.710 -20.920 ;
        RECT 120.110 -21.110 120.570 -20.920 ;
        RECT 117.260 -21.340 120.570 -21.110 ;
        RECT 117.260 -21.430 117.710 -21.340 ;
        RECT 120.110 -21.420 120.570 -21.340 ;
        RECT 124.060 -20.690 124.520 -20.610 ;
        RECT 126.920 -20.690 127.370 -20.600 ;
        RECT 124.060 -20.920 127.370 -20.690 ;
        RECT 124.060 -21.110 124.520 -20.920 ;
        RECT 126.920 -21.110 127.370 -20.920 ;
        RECT 124.060 -21.340 127.370 -21.110 ;
        RECT 124.060 -21.420 124.520 -21.340 ;
        RECT 126.920 -21.430 127.370 -21.340 ;
        RECT 130.760 -20.690 131.210 -20.600 ;
        RECT 133.610 -20.690 134.070 -20.610 ;
        RECT 130.760 -20.920 134.070 -20.690 ;
        RECT 130.760 -21.110 131.210 -20.920 ;
        RECT 133.610 -21.110 134.070 -20.920 ;
        RECT 130.760 -21.340 134.070 -21.110 ;
        RECT 130.760 -21.430 131.210 -21.340 ;
        RECT 133.610 -21.420 134.070 -21.340 ;
        RECT 137.560 -20.690 138.020 -20.610 ;
        RECT 140.420 -20.690 140.870 -20.600 ;
        RECT 137.560 -20.920 140.870 -20.690 ;
        RECT 137.560 -21.110 138.020 -20.920 ;
        RECT 140.420 -21.110 140.870 -20.920 ;
        RECT 137.560 -21.340 140.870 -21.110 ;
        RECT 137.560 -21.420 138.020 -21.340 ;
        RECT 140.420 -21.430 140.870 -21.340 ;
        RECT 144.260 -20.690 144.710 -20.600 ;
        RECT 147.110 -20.690 147.570 -20.610 ;
        RECT 144.260 -20.920 147.570 -20.690 ;
        RECT 144.260 -21.110 144.710 -20.920 ;
        RECT 147.110 -21.110 147.570 -20.920 ;
        RECT 144.260 -21.340 147.570 -21.110 ;
        RECT 144.260 -21.430 144.710 -21.340 ;
        RECT 147.110 -21.420 147.570 -21.340 ;
        RECT 151.060 -20.690 151.520 -20.610 ;
        RECT 153.920 -20.690 154.370 -20.600 ;
        RECT 151.060 -20.920 154.370 -20.690 ;
        RECT 151.060 -21.110 151.520 -20.920 ;
        RECT 153.920 -21.110 154.370 -20.920 ;
        RECT 151.060 -21.340 154.370 -21.110 ;
        RECT 151.060 -21.420 151.520 -21.340 ;
        RECT 153.920 -21.430 154.370 -21.340 ;
        RECT 157.760 -20.690 158.210 -20.600 ;
        RECT 160.610 -20.690 161.070 -20.610 ;
        RECT 157.760 -20.920 161.070 -20.690 ;
        RECT 157.760 -21.110 158.210 -20.920 ;
        RECT 160.610 -21.110 161.070 -20.920 ;
        RECT 157.760 -21.340 161.070 -21.110 ;
        RECT 157.760 -21.430 158.210 -21.340 ;
        RECT 160.610 -21.420 161.070 -21.340 ;
        RECT 164.560 -20.690 165.020 -20.610 ;
        RECT 167.420 -20.690 167.870 -20.600 ;
        RECT 164.560 -20.920 167.870 -20.690 ;
        RECT 164.560 -21.110 165.020 -20.920 ;
        RECT 167.420 -21.110 167.870 -20.920 ;
        RECT 164.560 -21.340 167.870 -21.110 ;
        RECT 164.560 -21.420 165.020 -21.340 ;
        RECT 167.420 -21.430 167.870 -21.340 ;
        RECT 171.260 -20.690 171.710 -20.600 ;
        RECT 174.110 -20.690 174.570 -20.610 ;
        RECT 171.260 -20.920 174.570 -20.690 ;
        RECT 171.260 -21.110 171.710 -20.920 ;
        RECT 174.110 -21.110 174.570 -20.920 ;
        RECT 171.260 -21.340 174.570 -21.110 ;
        RECT 171.260 -21.430 171.710 -21.340 ;
        RECT 174.110 -21.420 174.570 -21.340 ;
        RECT 178.060 -20.690 178.520 -20.610 ;
        RECT 180.920 -20.690 181.370 -20.600 ;
        RECT 178.060 -20.920 181.370 -20.690 ;
        RECT 178.060 -21.110 178.520 -20.920 ;
        RECT 180.920 -21.110 181.370 -20.920 ;
        RECT 178.060 -21.340 181.370 -21.110 ;
        RECT 178.060 -21.420 178.520 -21.340 ;
        RECT 180.920 -21.430 181.370 -21.340 ;
        RECT 184.760 -20.690 185.210 -20.600 ;
        RECT 187.610 -20.690 188.070 -20.610 ;
        RECT 184.760 -20.920 188.070 -20.690 ;
        RECT 184.760 -21.110 185.210 -20.920 ;
        RECT 187.610 -21.110 188.070 -20.920 ;
        RECT 184.760 -21.340 188.070 -21.110 ;
        RECT 184.760 -21.430 185.210 -21.340 ;
        RECT 187.610 -21.420 188.070 -21.340 ;
        RECT 191.560 -20.690 192.020 -20.610 ;
        RECT 194.420 -20.690 194.870 -20.600 ;
        RECT 191.560 -20.920 194.870 -20.690 ;
        RECT 191.560 -21.110 192.020 -20.920 ;
        RECT 194.420 -21.110 194.870 -20.920 ;
        RECT 191.560 -21.340 194.870 -21.110 ;
        RECT 191.560 -21.420 192.020 -21.340 ;
        RECT 194.420 -21.430 194.870 -21.340 ;
        RECT 198.260 -20.690 198.710 -20.600 ;
        RECT 201.110 -20.690 201.570 -20.610 ;
        RECT 198.260 -20.920 201.570 -20.690 ;
        RECT 198.260 -21.110 198.710 -20.920 ;
        RECT 201.110 -21.110 201.570 -20.920 ;
        RECT 198.260 -21.340 201.570 -21.110 ;
        RECT 198.260 -21.430 198.710 -21.340 ;
        RECT 201.110 -21.420 201.570 -21.340 ;
        RECT 205.060 -20.690 205.520 -20.610 ;
        RECT 207.920 -20.690 208.370 -20.600 ;
        RECT 205.060 -20.920 208.370 -20.690 ;
        RECT 205.060 -21.110 205.520 -20.920 ;
        RECT 207.920 -21.110 208.370 -20.920 ;
        RECT 205.060 -21.340 208.370 -21.110 ;
        RECT 205.060 -21.420 205.520 -21.340 ;
        RECT 207.920 -21.430 208.370 -21.340 ;
        RECT 211.760 -20.690 212.210 -20.600 ;
        RECT 214.610 -20.690 215.070 -20.610 ;
        RECT 211.760 -20.920 215.070 -20.690 ;
        RECT 211.760 -21.110 212.210 -20.920 ;
        RECT 214.610 -21.110 215.070 -20.920 ;
        RECT 211.760 -21.340 215.070 -21.110 ;
        RECT 211.760 -21.430 212.210 -21.340 ;
        RECT 214.610 -21.420 215.070 -21.340 ;
        RECT 9.260 -24.300 9.710 -24.210 ;
        RECT 12.110 -24.300 12.570 -24.220 ;
        RECT 9.260 -24.530 12.570 -24.300 ;
        RECT 9.260 -24.720 9.710 -24.530 ;
        RECT 12.110 -24.720 12.570 -24.530 ;
        RECT 9.260 -24.950 12.570 -24.720 ;
        RECT 9.260 -25.040 9.710 -24.950 ;
        RECT 12.110 -25.030 12.570 -24.950 ;
        RECT 16.060 -24.300 16.520 -24.220 ;
        RECT 18.920 -24.300 19.370 -24.210 ;
        RECT 16.060 -24.530 19.370 -24.300 ;
        RECT 16.060 -24.720 16.520 -24.530 ;
        RECT 18.920 -24.720 19.370 -24.530 ;
        RECT 16.060 -24.950 19.370 -24.720 ;
        RECT 16.060 -25.030 16.520 -24.950 ;
        RECT 18.920 -25.040 19.370 -24.950 ;
        RECT 22.760 -24.300 23.210 -24.210 ;
        RECT 25.610 -24.300 26.070 -24.220 ;
        RECT 22.760 -24.530 26.070 -24.300 ;
        RECT 22.760 -24.720 23.210 -24.530 ;
        RECT 25.610 -24.720 26.070 -24.530 ;
        RECT 22.760 -24.950 26.070 -24.720 ;
        RECT 22.760 -25.040 23.210 -24.950 ;
        RECT 25.610 -25.030 26.070 -24.950 ;
        RECT 29.560 -24.300 30.020 -24.220 ;
        RECT 32.420 -24.300 32.870 -24.210 ;
        RECT 29.560 -24.530 32.870 -24.300 ;
        RECT 29.560 -24.720 30.020 -24.530 ;
        RECT 32.420 -24.720 32.870 -24.530 ;
        RECT 29.560 -24.950 32.870 -24.720 ;
        RECT 29.560 -25.030 30.020 -24.950 ;
        RECT 32.420 -25.040 32.870 -24.950 ;
        RECT 36.260 -24.300 36.710 -24.210 ;
        RECT 39.110 -24.300 39.570 -24.220 ;
        RECT 36.260 -24.530 39.570 -24.300 ;
        RECT 36.260 -24.720 36.710 -24.530 ;
        RECT 39.110 -24.720 39.570 -24.530 ;
        RECT 36.260 -24.950 39.570 -24.720 ;
        RECT 36.260 -25.040 36.710 -24.950 ;
        RECT 39.110 -25.030 39.570 -24.950 ;
        RECT 43.060 -24.300 43.520 -24.220 ;
        RECT 45.920 -24.300 46.370 -24.210 ;
        RECT 43.060 -24.530 46.370 -24.300 ;
        RECT 43.060 -24.720 43.520 -24.530 ;
        RECT 45.920 -24.720 46.370 -24.530 ;
        RECT 43.060 -24.950 46.370 -24.720 ;
        RECT 43.060 -25.030 43.520 -24.950 ;
        RECT 45.920 -25.040 46.370 -24.950 ;
        RECT 49.760 -24.300 50.210 -24.210 ;
        RECT 52.610 -24.300 53.070 -24.220 ;
        RECT 49.760 -24.530 53.070 -24.300 ;
        RECT 49.760 -24.720 50.210 -24.530 ;
        RECT 52.610 -24.720 53.070 -24.530 ;
        RECT 49.760 -24.950 53.070 -24.720 ;
        RECT 49.760 -25.040 50.210 -24.950 ;
        RECT 52.610 -25.030 53.070 -24.950 ;
        RECT 56.560 -24.300 57.020 -24.220 ;
        RECT 59.420 -24.300 59.870 -24.210 ;
        RECT 56.560 -24.530 59.870 -24.300 ;
        RECT 56.560 -24.720 57.020 -24.530 ;
        RECT 59.420 -24.720 59.870 -24.530 ;
        RECT 56.560 -24.950 59.870 -24.720 ;
        RECT 56.560 -25.030 57.020 -24.950 ;
        RECT 59.420 -25.040 59.870 -24.950 ;
        RECT 63.260 -24.300 63.710 -24.210 ;
        RECT 66.110 -24.300 66.570 -24.220 ;
        RECT 63.260 -24.530 66.570 -24.300 ;
        RECT 63.260 -24.720 63.710 -24.530 ;
        RECT 66.110 -24.720 66.570 -24.530 ;
        RECT 63.260 -24.950 66.570 -24.720 ;
        RECT 63.260 -25.040 63.710 -24.950 ;
        RECT 66.110 -25.030 66.570 -24.950 ;
        RECT 70.060 -24.300 70.520 -24.220 ;
        RECT 72.920 -24.300 73.370 -24.210 ;
        RECT 70.060 -24.530 73.370 -24.300 ;
        RECT 70.060 -24.720 70.520 -24.530 ;
        RECT 72.920 -24.720 73.370 -24.530 ;
        RECT 70.060 -24.950 73.370 -24.720 ;
        RECT 70.060 -25.030 70.520 -24.950 ;
        RECT 72.920 -25.040 73.370 -24.950 ;
        RECT 76.760 -24.300 77.210 -24.210 ;
        RECT 79.610 -24.300 80.070 -24.220 ;
        RECT 76.760 -24.530 80.070 -24.300 ;
        RECT 76.760 -24.720 77.210 -24.530 ;
        RECT 79.610 -24.720 80.070 -24.530 ;
        RECT 76.760 -24.950 80.070 -24.720 ;
        RECT 76.760 -25.040 77.210 -24.950 ;
        RECT 79.610 -25.030 80.070 -24.950 ;
        RECT 83.560 -24.300 84.020 -24.220 ;
        RECT 86.420 -24.300 86.870 -24.210 ;
        RECT 83.560 -24.530 86.870 -24.300 ;
        RECT 83.560 -24.720 84.020 -24.530 ;
        RECT 86.420 -24.720 86.870 -24.530 ;
        RECT 83.560 -24.950 86.870 -24.720 ;
        RECT 83.560 -25.030 84.020 -24.950 ;
        RECT 86.420 -25.040 86.870 -24.950 ;
        RECT 90.260 -24.300 90.710 -24.210 ;
        RECT 93.110 -24.300 93.570 -24.220 ;
        RECT 90.260 -24.530 93.570 -24.300 ;
        RECT 90.260 -24.720 90.710 -24.530 ;
        RECT 93.110 -24.720 93.570 -24.530 ;
        RECT 90.260 -24.950 93.570 -24.720 ;
        RECT 90.260 -25.040 90.710 -24.950 ;
        RECT 93.110 -25.030 93.570 -24.950 ;
        RECT 97.060 -24.300 97.520 -24.220 ;
        RECT 99.920 -24.300 100.370 -24.210 ;
        RECT 97.060 -24.530 100.370 -24.300 ;
        RECT 97.060 -24.720 97.520 -24.530 ;
        RECT 99.920 -24.720 100.370 -24.530 ;
        RECT 97.060 -24.950 100.370 -24.720 ;
        RECT 97.060 -25.030 97.520 -24.950 ;
        RECT 99.920 -25.040 100.370 -24.950 ;
        RECT 103.760 -24.300 104.210 -24.210 ;
        RECT 106.610 -24.300 107.070 -24.220 ;
        RECT 103.760 -24.530 107.070 -24.300 ;
        RECT 103.760 -24.720 104.210 -24.530 ;
        RECT 106.610 -24.720 107.070 -24.530 ;
        RECT 103.760 -24.950 107.070 -24.720 ;
        RECT 103.760 -25.040 104.210 -24.950 ;
        RECT 106.610 -25.030 107.070 -24.950 ;
        RECT 110.560 -24.300 111.020 -24.220 ;
        RECT 113.420 -24.300 113.870 -24.210 ;
        RECT 110.560 -24.530 113.870 -24.300 ;
        RECT 110.560 -24.720 111.020 -24.530 ;
        RECT 113.420 -24.720 113.870 -24.530 ;
        RECT 110.560 -24.950 113.870 -24.720 ;
        RECT 110.560 -25.030 111.020 -24.950 ;
        RECT 113.420 -25.040 113.870 -24.950 ;
        RECT 117.260 -24.300 117.710 -24.210 ;
        RECT 120.110 -24.300 120.570 -24.220 ;
        RECT 117.260 -24.530 120.570 -24.300 ;
        RECT 117.260 -24.720 117.710 -24.530 ;
        RECT 120.110 -24.720 120.570 -24.530 ;
        RECT 117.260 -24.950 120.570 -24.720 ;
        RECT 117.260 -25.040 117.710 -24.950 ;
        RECT 120.110 -25.030 120.570 -24.950 ;
        RECT 124.060 -24.300 124.520 -24.220 ;
        RECT 126.920 -24.300 127.370 -24.210 ;
        RECT 124.060 -24.530 127.370 -24.300 ;
        RECT 124.060 -24.720 124.520 -24.530 ;
        RECT 126.920 -24.720 127.370 -24.530 ;
        RECT 124.060 -24.950 127.370 -24.720 ;
        RECT 124.060 -25.030 124.520 -24.950 ;
        RECT 126.920 -25.040 127.370 -24.950 ;
        RECT 130.760 -24.300 131.210 -24.210 ;
        RECT 133.610 -24.300 134.070 -24.220 ;
        RECT 130.760 -24.530 134.070 -24.300 ;
        RECT 130.760 -24.720 131.210 -24.530 ;
        RECT 133.610 -24.720 134.070 -24.530 ;
        RECT 130.760 -24.950 134.070 -24.720 ;
        RECT 130.760 -25.040 131.210 -24.950 ;
        RECT 133.610 -25.030 134.070 -24.950 ;
        RECT 137.560 -24.300 138.020 -24.220 ;
        RECT 140.420 -24.300 140.870 -24.210 ;
        RECT 137.560 -24.530 140.870 -24.300 ;
        RECT 137.560 -24.720 138.020 -24.530 ;
        RECT 140.420 -24.720 140.870 -24.530 ;
        RECT 137.560 -24.950 140.870 -24.720 ;
        RECT 137.560 -25.030 138.020 -24.950 ;
        RECT 140.420 -25.040 140.870 -24.950 ;
        RECT 144.260 -24.300 144.710 -24.210 ;
        RECT 147.110 -24.300 147.570 -24.220 ;
        RECT 144.260 -24.530 147.570 -24.300 ;
        RECT 144.260 -24.720 144.710 -24.530 ;
        RECT 147.110 -24.720 147.570 -24.530 ;
        RECT 144.260 -24.950 147.570 -24.720 ;
        RECT 144.260 -25.040 144.710 -24.950 ;
        RECT 147.110 -25.030 147.570 -24.950 ;
        RECT 151.060 -24.300 151.520 -24.220 ;
        RECT 153.920 -24.300 154.370 -24.210 ;
        RECT 151.060 -24.530 154.370 -24.300 ;
        RECT 151.060 -24.720 151.520 -24.530 ;
        RECT 153.920 -24.720 154.370 -24.530 ;
        RECT 151.060 -24.950 154.370 -24.720 ;
        RECT 151.060 -25.030 151.520 -24.950 ;
        RECT 153.920 -25.040 154.370 -24.950 ;
        RECT 157.760 -24.300 158.210 -24.210 ;
        RECT 160.610 -24.300 161.070 -24.220 ;
        RECT 157.760 -24.530 161.070 -24.300 ;
        RECT 157.760 -24.720 158.210 -24.530 ;
        RECT 160.610 -24.720 161.070 -24.530 ;
        RECT 157.760 -24.950 161.070 -24.720 ;
        RECT 157.760 -25.040 158.210 -24.950 ;
        RECT 160.610 -25.030 161.070 -24.950 ;
        RECT 164.560 -24.300 165.020 -24.220 ;
        RECT 167.420 -24.300 167.870 -24.210 ;
        RECT 164.560 -24.530 167.870 -24.300 ;
        RECT 164.560 -24.720 165.020 -24.530 ;
        RECT 167.420 -24.720 167.870 -24.530 ;
        RECT 164.560 -24.950 167.870 -24.720 ;
        RECT 164.560 -25.030 165.020 -24.950 ;
        RECT 167.420 -25.040 167.870 -24.950 ;
        RECT 171.260 -24.300 171.710 -24.210 ;
        RECT 174.110 -24.300 174.570 -24.220 ;
        RECT 171.260 -24.530 174.570 -24.300 ;
        RECT 171.260 -24.720 171.710 -24.530 ;
        RECT 174.110 -24.720 174.570 -24.530 ;
        RECT 171.260 -24.950 174.570 -24.720 ;
        RECT 171.260 -25.040 171.710 -24.950 ;
        RECT 174.110 -25.030 174.570 -24.950 ;
        RECT 178.060 -24.300 178.520 -24.220 ;
        RECT 180.920 -24.300 181.370 -24.210 ;
        RECT 178.060 -24.530 181.370 -24.300 ;
        RECT 178.060 -24.720 178.520 -24.530 ;
        RECT 180.920 -24.720 181.370 -24.530 ;
        RECT 178.060 -24.950 181.370 -24.720 ;
        RECT 178.060 -25.030 178.520 -24.950 ;
        RECT 180.920 -25.040 181.370 -24.950 ;
        RECT 184.760 -24.300 185.210 -24.210 ;
        RECT 187.610 -24.300 188.070 -24.220 ;
        RECT 184.760 -24.530 188.070 -24.300 ;
        RECT 184.760 -24.720 185.210 -24.530 ;
        RECT 187.610 -24.720 188.070 -24.530 ;
        RECT 184.760 -24.950 188.070 -24.720 ;
        RECT 184.760 -25.040 185.210 -24.950 ;
        RECT 187.610 -25.030 188.070 -24.950 ;
        RECT 191.560 -24.300 192.020 -24.220 ;
        RECT 194.420 -24.300 194.870 -24.210 ;
        RECT 191.560 -24.530 194.870 -24.300 ;
        RECT 191.560 -24.720 192.020 -24.530 ;
        RECT 194.420 -24.720 194.870 -24.530 ;
        RECT 191.560 -24.950 194.870 -24.720 ;
        RECT 191.560 -25.030 192.020 -24.950 ;
        RECT 194.420 -25.040 194.870 -24.950 ;
        RECT 198.260 -24.300 198.710 -24.210 ;
        RECT 201.110 -24.300 201.570 -24.220 ;
        RECT 198.260 -24.530 201.570 -24.300 ;
        RECT 198.260 -24.720 198.710 -24.530 ;
        RECT 201.110 -24.720 201.570 -24.530 ;
        RECT 198.260 -24.950 201.570 -24.720 ;
        RECT 198.260 -25.040 198.710 -24.950 ;
        RECT 201.110 -25.030 201.570 -24.950 ;
        RECT 205.060 -24.300 205.520 -24.220 ;
        RECT 207.920 -24.300 208.370 -24.210 ;
        RECT 205.060 -24.530 208.370 -24.300 ;
        RECT 205.060 -24.720 205.520 -24.530 ;
        RECT 207.920 -24.720 208.370 -24.530 ;
        RECT 205.060 -24.950 208.370 -24.720 ;
        RECT 205.060 -25.030 205.520 -24.950 ;
        RECT 207.920 -25.040 208.370 -24.950 ;
        RECT 211.760 -24.300 212.210 -24.210 ;
        RECT 214.610 -24.300 215.070 -24.220 ;
        RECT 211.760 -24.530 215.070 -24.300 ;
        RECT 211.760 -24.720 212.210 -24.530 ;
        RECT 214.610 -24.720 215.070 -24.530 ;
        RECT 211.760 -24.950 215.070 -24.720 ;
        RECT 211.760 -25.040 212.210 -24.950 ;
        RECT 214.610 -25.030 215.070 -24.950 ;
        RECT 9.260 -27.910 9.710 -27.820 ;
        RECT 12.110 -27.910 12.570 -27.830 ;
        RECT 9.260 -28.140 12.570 -27.910 ;
        RECT 9.260 -28.330 9.710 -28.140 ;
        RECT 12.110 -28.330 12.570 -28.140 ;
        RECT 9.260 -28.560 12.570 -28.330 ;
        RECT 9.260 -28.650 9.710 -28.560 ;
        RECT 12.110 -28.640 12.570 -28.560 ;
        RECT 16.060 -27.910 16.520 -27.830 ;
        RECT 18.920 -27.910 19.370 -27.820 ;
        RECT 16.060 -28.140 19.370 -27.910 ;
        RECT 16.060 -28.330 16.520 -28.140 ;
        RECT 18.920 -28.330 19.370 -28.140 ;
        RECT 16.060 -28.560 19.370 -28.330 ;
        RECT 16.060 -28.640 16.520 -28.560 ;
        RECT 18.920 -28.650 19.370 -28.560 ;
        RECT 22.760 -27.910 23.210 -27.820 ;
        RECT 25.610 -27.910 26.070 -27.830 ;
        RECT 22.760 -28.140 26.070 -27.910 ;
        RECT 22.760 -28.330 23.210 -28.140 ;
        RECT 25.610 -28.330 26.070 -28.140 ;
        RECT 22.760 -28.560 26.070 -28.330 ;
        RECT 22.760 -28.650 23.210 -28.560 ;
        RECT 25.610 -28.640 26.070 -28.560 ;
        RECT 29.560 -27.910 30.020 -27.830 ;
        RECT 32.420 -27.910 32.870 -27.820 ;
        RECT 29.560 -28.140 32.870 -27.910 ;
        RECT 29.560 -28.330 30.020 -28.140 ;
        RECT 32.420 -28.330 32.870 -28.140 ;
        RECT 29.560 -28.560 32.870 -28.330 ;
        RECT 29.560 -28.640 30.020 -28.560 ;
        RECT 32.420 -28.650 32.870 -28.560 ;
        RECT 36.260 -27.910 36.710 -27.820 ;
        RECT 39.110 -27.910 39.570 -27.830 ;
        RECT 36.260 -28.140 39.570 -27.910 ;
        RECT 36.260 -28.330 36.710 -28.140 ;
        RECT 39.110 -28.330 39.570 -28.140 ;
        RECT 36.260 -28.560 39.570 -28.330 ;
        RECT 36.260 -28.650 36.710 -28.560 ;
        RECT 39.110 -28.640 39.570 -28.560 ;
        RECT 43.060 -27.910 43.520 -27.830 ;
        RECT 45.920 -27.910 46.370 -27.820 ;
        RECT 43.060 -28.140 46.370 -27.910 ;
        RECT 43.060 -28.330 43.520 -28.140 ;
        RECT 45.920 -28.330 46.370 -28.140 ;
        RECT 43.060 -28.560 46.370 -28.330 ;
        RECT 43.060 -28.640 43.520 -28.560 ;
        RECT 45.920 -28.650 46.370 -28.560 ;
        RECT 49.760 -27.910 50.210 -27.820 ;
        RECT 52.610 -27.910 53.070 -27.830 ;
        RECT 49.760 -28.140 53.070 -27.910 ;
        RECT 49.760 -28.330 50.210 -28.140 ;
        RECT 52.610 -28.330 53.070 -28.140 ;
        RECT 49.760 -28.560 53.070 -28.330 ;
        RECT 49.760 -28.650 50.210 -28.560 ;
        RECT 52.610 -28.640 53.070 -28.560 ;
        RECT 56.560 -27.910 57.020 -27.830 ;
        RECT 59.420 -27.910 59.870 -27.820 ;
        RECT 56.560 -28.140 59.870 -27.910 ;
        RECT 56.560 -28.330 57.020 -28.140 ;
        RECT 59.420 -28.330 59.870 -28.140 ;
        RECT 56.560 -28.560 59.870 -28.330 ;
        RECT 56.560 -28.640 57.020 -28.560 ;
        RECT 59.420 -28.650 59.870 -28.560 ;
        RECT 63.260 -27.910 63.710 -27.820 ;
        RECT 66.110 -27.910 66.570 -27.830 ;
        RECT 63.260 -28.140 66.570 -27.910 ;
        RECT 63.260 -28.330 63.710 -28.140 ;
        RECT 66.110 -28.330 66.570 -28.140 ;
        RECT 63.260 -28.560 66.570 -28.330 ;
        RECT 63.260 -28.650 63.710 -28.560 ;
        RECT 66.110 -28.640 66.570 -28.560 ;
        RECT 70.060 -27.910 70.520 -27.830 ;
        RECT 72.920 -27.910 73.370 -27.820 ;
        RECT 70.060 -28.140 73.370 -27.910 ;
        RECT 70.060 -28.330 70.520 -28.140 ;
        RECT 72.920 -28.330 73.370 -28.140 ;
        RECT 70.060 -28.560 73.370 -28.330 ;
        RECT 70.060 -28.640 70.520 -28.560 ;
        RECT 72.920 -28.650 73.370 -28.560 ;
        RECT 76.760 -27.910 77.210 -27.820 ;
        RECT 79.610 -27.910 80.070 -27.830 ;
        RECT 76.760 -28.140 80.070 -27.910 ;
        RECT 76.760 -28.330 77.210 -28.140 ;
        RECT 79.610 -28.330 80.070 -28.140 ;
        RECT 76.760 -28.560 80.070 -28.330 ;
        RECT 76.760 -28.650 77.210 -28.560 ;
        RECT 79.610 -28.640 80.070 -28.560 ;
        RECT 83.560 -27.910 84.020 -27.830 ;
        RECT 86.420 -27.910 86.870 -27.820 ;
        RECT 83.560 -28.140 86.870 -27.910 ;
        RECT 83.560 -28.330 84.020 -28.140 ;
        RECT 86.420 -28.330 86.870 -28.140 ;
        RECT 83.560 -28.560 86.870 -28.330 ;
        RECT 83.560 -28.640 84.020 -28.560 ;
        RECT 86.420 -28.650 86.870 -28.560 ;
        RECT 90.260 -27.910 90.710 -27.820 ;
        RECT 93.110 -27.910 93.570 -27.830 ;
        RECT 90.260 -28.140 93.570 -27.910 ;
        RECT 90.260 -28.330 90.710 -28.140 ;
        RECT 93.110 -28.330 93.570 -28.140 ;
        RECT 90.260 -28.560 93.570 -28.330 ;
        RECT 90.260 -28.650 90.710 -28.560 ;
        RECT 93.110 -28.640 93.570 -28.560 ;
        RECT 97.060 -27.910 97.520 -27.830 ;
        RECT 99.920 -27.910 100.370 -27.820 ;
        RECT 97.060 -28.140 100.370 -27.910 ;
        RECT 97.060 -28.330 97.520 -28.140 ;
        RECT 99.920 -28.330 100.370 -28.140 ;
        RECT 97.060 -28.560 100.370 -28.330 ;
        RECT 97.060 -28.640 97.520 -28.560 ;
        RECT 99.920 -28.650 100.370 -28.560 ;
        RECT 103.760 -27.910 104.210 -27.820 ;
        RECT 106.610 -27.910 107.070 -27.830 ;
        RECT 103.760 -28.140 107.070 -27.910 ;
        RECT 103.760 -28.330 104.210 -28.140 ;
        RECT 106.610 -28.330 107.070 -28.140 ;
        RECT 103.760 -28.560 107.070 -28.330 ;
        RECT 103.760 -28.650 104.210 -28.560 ;
        RECT 106.610 -28.640 107.070 -28.560 ;
        RECT 110.560 -27.910 111.020 -27.830 ;
        RECT 113.420 -27.910 113.870 -27.820 ;
        RECT 110.560 -28.140 113.870 -27.910 ;
        RECT 110.560 -28.330 111.020 -28.140 ;
        RECT 113.420 -28.330 113.870 -28.140 ;
        RECT 110.560 -28.560 113.870 -28.330 ;
        RECT 110.560 -28.640 111.020 -28.560 ;
        RECT 113.420 -28.650 113.870 -28.560 ;
        RECT 117.260 -27.910 117.710 -27.820 ;
        RECT 120.110 -27.910 120.570 -27.830 ;
        RECT 117.260 -28.140 120.570 -27.910 ;
        RECT 117.260 -28.330 117.710 -28.140 ;
        RECT 120.110 -28.330 120.570 -28.140 ;
        RECT 117.260 -28.560 120.570 -28.330 ;
        RECT 117.260 -28.650 117.710 -28.560 ;
        RECT 120.110 -28.640 120.570 -28.560 ;
        RECT 124.060 -27.910 124.520 -27.830 ;
        RECT 126.920 -27.910 127.370 -27.820 ;
        RECT 124.060 -28.140 127.370 -27.910 ;
        RECT 124.060 -28.330 124.520 -28.140 ;
        RECT 126.920 -28.330 127.370 -28.140 ;
        RECT 124.060 -28.560 127.370 -28.330 ;
        RECT 124.060 -28.640 124.520 -28.560 ;
        RECT 126.920 -28.650 127.370 -28.560 ;
        RECT 130.760 -27.910 131.210 -27.820 ;
        RECT 133.610 -27.910 134.070 -27.830 ;
        RECT 130.760 -28.140 134.070 -27.910 ;
        RECT 130.760 -28.330 131.210 -28.140 ;
        RECT 133.610 -28.330 134.070 -28.140 ;
        RECT 130.760 -28.560 134.070 -28.330 ;
        RECT 130.760 -28.650 131.210 -28.560 ;
        RECT 133.610 -28.640 134.070 -28.560 ;
        RECT 137.560 -27.910 138.020 -27.830 ;
        RECT 140.420 -27.910 140.870 -27.820 ;
        RECT 137.560 -28.140 140.870 -27.910 ;
        RECT 137.560 -28.330 138.020 -28.140 ;
        RECT 140.420 -28.330 140.870 -28.140 ;
        RECT 137.560 -28.560 140.870 -28.330 ;
        RECT 137.560 -28.640 138.020 -28.560 ;
        RECT 140.420 -28.650 140.870 -28.560 ;
        RECT 144.260 -27.910 144.710 -27.820 ;
        RECT 147.110 -27.910 147.570 -27.830 ;
        RECT 144.260 -28.140 147.570 -27.910 ;
        RECT 144.260 -28.330 144.710 -28.140 ;
        RECT 147.110 -28.330 147.570 -28.140 ;
        RECT 144.260 -28.560 147.570 -28.330 ;
        RECT 144.260 -28.650 144.710 -28.560 ;
        RECT 147.110 -28.640 147.570 -28.560 ;
        RECT 151.060 -27.910 151.520 -27.830 ;
        RECT 153.920 -27.910 154.370 -27.820 ;
        RECT 151.060 -28.140 154.370 -27.910 ;
        RECT 151.060 -28.330 151.520 -28.140 ;
        RECT 153.920 -28.330 154.370 -28.140 ;
        RECT 151.060 -28.560 154.370 -28.330 ;
        RECT 151.060 -28.640 151.520 -28.560 ;
        RECT 153.920 -28.650 154.370 -28.560 ;
        RECT 157.760 -27.910 158.210 -27.820 ;
        RECT 160.610 -27.910 161.070 -27.830 ;
        RECT 157.760 -28.140 161.070 -27.910 ;
        RECT 157.760 -28.330 158.210 -28.140 ;
        RECT 160.610 -28.330 161.070 -28.140 ;
        RECT 157.760 -28.560 161.070 -28.330 ;
        RECT 157.760 -28.650 158.210 -28.560 ;
        RECT 160.610 -28.640 161.070 -28.560 ;
        RECT 164.560 -27.910 165.020 -27.830 ;
        RECT 167.420 -27.910 167.870 -27.820 ;
        RECT 164.560 -28.140 167.870 -27.910 ;
        RECT 164.560 -28.330 165.020 -28.140 ;
        RECT 167.420 -28.330 167.870 -28.140 ;
        RECT 164.560 -28.560 167.870 -28.330 ;
        RECT 164.560 -28.640 165.020 -28.560 ;
        RECT 167.420 -28.650 167.870 -28.560 ;
        RECT 171.260 -27.910 171.710 -27.820 ;
        RECT 174.110 -27.910 174.570 -27.830 ;
        RECT 171.260 -28.140 174.570 -27.910 ;
        RECT 171.260 -28.330 171.710 -28.140 ;
        RECT 174.110 -28.330 174.570 -28.140 ;
        RECT 171.260 -28.560 174.570 -28.330 ;
        RECT 171.260 -28.650 171.710 -28.560 ;
        RECT 174.110 -28.640 174.570 -28.560 ;
        RECT 178.060 -27.910 178.520 -27.830 ;
        RECT 180.920 -27.910 181.370 -27.820 ;
        RECT 178.060 -28.140 181.370 -27.910 ;
        RECT 178.060 -28.330 178.520 -28.140 ;
        RECT 180.920 -28.330 181.370 -28.140 ;
        RECT 178.060 -28.560 181.370 -28.330 ;
        RECT 178.060 -28.640 178.520 -28.560 ;
        RECT 180.920 -28.650 181.370 -28.560 ;
        RECT 184.760 -27.910 185.210 -27.820 ;
        RECT 187.610 -27.910 188.070 -27.830 ;
        RECT 184.760 -28.140 188.070 -27.910 ;
        RECT 184.760 -28.330 185.210 -28.140 ;
        RECT 187.610 -28.330 188.070 -28.140 ;
        RECT 184.760 -28.560 188.070 -28.330 ;
        RECT 184.760 -28.650 185.210 -28.560 ;
        RECT 187.610 -28.640 188.070 -28.560 ;
        RECT 191.560 -27.910 192.020 -27.830 ;
        RECT 194.420 -27.910 194.870 -27.820 ;
        RECT 191.560 -28.140 194.870 -27.910 ;
        RECT 191.560 -28.330 192.020 -28.140 ;
        RECT 194.420 -28.330 194.870 -28.140 ;
        RECT 191.560 -28.560 194.870 -28.330 ;
        RECT 191.560 -28.640 192.020 -28.560 ;
        RECT 194.420 -28.650 194.870 -28.560 ;
        RECT 198.260 -27.910 198.710 -27.820 ;
        RECT 201.110 -27.910 201.570 -27.830 ;
        RECT 198.260 -28.140 201.570 -27.910 ;
        RECT 198.260 -28.330 198.710 -28.140 ;
        RECT 201.110 -28.330 201.570 -28.140 ;
        RECT 198.260 -28.560 201.570 -28.330 ;
        RECT 198.260 -28.650 198.710 -28.560 ;
        RECT 201.110 -28.640 201.570 -28.560 ;
        RECT 205.060 -27.910 205.520 -27.830 ;
        RECT 207.920 -27.910 208.370 -27.820 ;
        RECT 205.060 -28.140 208.370 -27.910 ;
        RECT 205.060 -28.330 205.520 -28.140 ;
        RECT 207.920 -28.330 208.370 -28.140 ;
        RECT 205.060 -28.560 208.370 -28.330 ;
        RECT 205.060 -28.640 205.520 -28.560 ;
        RECT 207.920 -28.650 208.370 -28.560 ;
        RECT 211.760 -27.910 212.210 -27.820 ;
        RECT 214.610 -27.910 215.070 -27.830 ;
        RECT 211.760 -28.140 215.070 -27.910 ;
        RECT 211.760 -28.330 212.210 -28.140 ;
        RECT 214.610 -28.330 215.070 -28.140 ;
        RECT 211.760 -28.560 215.070 -28.330 ;
        RECT 211.760 -28.650 212.210 -28.560 ;
        RECT 214.610 -28.640 215.070 -28.560 ;
        RECT 9.260 -31.520 9.710 -31.430 ;
        RECT 12.110 -31.520 12.570 -31.440 ;
        RECT 9.260 -31.750 12.570 -31.520 ;
        RECT 9.260 -31.940 9.710 -31.750 ;
        RECT 12.110 -31.940 12.570 -31.750 ;
        RECT 9.260 -32.170 12.570 -31.940 ;
        RECT 9.260 -32.260 9.710 -32.170 ;
        RECT 12.110 -32.250 12.570 -32.170 ;
        RECT 16.060 -31.520 16.520 -31.440 ;
        RECT 18.920 -31.520 19.370 -31.430 ;
        RECT 16.060 -31.750 19.370 -31.520 ;
        RECT 16.060 -31.940 16.520 -31.750 ;
        RECT 18.920 -31.940 19.370 -31.750 ;
        RECT 16.060 -32.170 19.370 -31.940 ;
        RECT 16.060 -32.250 16.520 -32.170 ;
        RECT 18.920 -32.260 19.370 -32.170 ;
        RECT 22.760 -31.520 23.210 -31.430 ;
        RECT 25.610 -31.520 26.070 -31.440 ;
        RECT 22.760 -31.750 26.070 -31.520 ;
        RECT 22.760 -31.940 23.210 -31.750 ;
        RECT 25.610 -31.940 26.070 -31.750 ;
        RECT 22.760 -32.170 26.070 -31.940 ;
        RECT 22.760 -32.260 23.210 -32.170 ;
        RECT 25.610 -32.250 26.070 -32.170 ;
        RECT 29.560 -31.520 30.020 -31.440 ;
        RECT 32.420 -31.520 32.870 -31.430 ;
        RECT 29.560 -31.750 32.870 -31.520 ;
        RECT 29.560 -31.940 30.020 -31.750 ;
        RECT 32.420 -31.940 32.870 -31.750 ;
        RECT 29.560 -32.170 32.870 -31.940 ;
        RECT 29.560 -32.250 30.020 -32.170 ;
        RECT 32.420 -32.260 32.870 -32.170 ;
        RECT 36.260 -31.520 36.710 -31.430 ;
        RECT 39.110 -31.520 39.570 -31.440 ;
        RECT 36.260 -31.750 39.570 -31.520 ;
        RECT 36.260 -31.940 36.710 -31.750 ;
        RECT 39.110 -31.940 39.570 -31.750 ;
        RECT 36.260 -32.170 39.570 -31.940 ;
        RECT 36.260 -32.260 36.710 -32.170 ;
        RECT 39.110 -32.250 39.570 -32.170 ;
        RECT 43.060 -31.520 43.520 -31.440 ;
        RECT 45.920 -31.520 46.370 -31.430 ;
        RECT 43.060 -31.750 46.370 -31.520 ;
        RECT 43.060 -31.940 43.520 -31.750 ;
        RECT 45.920 -31.940 46.370 -31.750 ;
        RECT 43.060 -32.170 46.370 -31.940 ;
        RECT 43.060 -32.250 43.520 -32.170 ;
        RECT 45.920 -32.260 46.370 -32.170 ;
        RECT 49.760 -31.520 50.210 -31.430 ;
        RECT 52.610 -31.520 53.070 -31.440 ;
        RECT 49.760 -31.750 53.070 -31.520 ;
        RECT 49.760 -31.940 50.210 -31.750 ;
        RECT 52.610 -31.940 53.070 -31.750 ;
        RECT 49.760 -32.170 53.070 -31.940 ;
        RECT 49.760 -32.260 50.210 -32.170 ;
        RECT 52.610 -32.250 53.070 -32.170 ;
        RECT 56.560 -31.520 57.020 -31.440 ;
        RECT 59.420 -31.520 59.870 -31.430 ;
        RECT 56.560 -31.750 59.870 -31.520 ;
        RECT 56.560 -31.940 57.020 -31.750 ;
        RECT 59.420 -31.940 59.870 -31.750 ;
        RECT 56.560 -32.170 59.870 -31.940 ;
        RECT 56.560 -32.250 57.020 -32.170 ;
        RECT 59.420 -32.260 59.870 -32.170 ;
        RECT 63.260 -31.520 63.710 -31.430 ;
        RECT 66.110 -31.520 66.570 -31.440 ;
        RECT 63.260 -31.750 66.570 -31.520 ;
        RECT 63.260 -31.940 63.710 -31.750 ;
        RECT 66.110 -31.940 66.570 -31.750 ;
        RECT 63.260 -32.170 66.570 -31.940 ;
        RECT 63.260 -32.260 63.710 -32.170 ;
        RECT 66.110 -32.250 66.570 -32.170 ;
        RECT 70.060 -31.520 70.520 -31.440 ;
        RECT 72.920 -31.520 73.370 -31.430 ;
        RECT 70.060 -31.750 73.370 -31.520 ;
        RECT 70.060 -31.940 70.520 -31.750 ;
        RECT 72.920 -31.940 73.370 -31.750 ;
        RECT 70.060 -32.170 73.370 -31.940 ;
        RECT 70.060 -32.250 70.520 -32.170 ;
        RECT 72.920 -32.260 73.370 -32.170 ;
        RECT 76.760 -31.520 77.210 -31.430 ;
        RECT 79.610 -31.520 80.070 -31.440 ;
        RECT 76.760 -31.750 80.070 -31.520 ;
        RECT 76.760 -31.940 77.210 -31.750 ;
        RECT 79.610 -31.940 80.070 -31.750 ;
        RECT 76.760 -32.170 80.070 -31.940 ;
        RECT 76.760 -32.260 77.210 -32.170 ;
        RECT 79.610 -32.250 80.070 -32.170 ;
        RECT 83.560 -31.520 84.020 -31.440 ;
        RECT 86.420 -31.520 86.870 -31.430 ;
        RECT 83.560 -31.750 86.870 -31.520 ;
        RECT 83.560 -31.940 84.020 -31.750 ;
        RECT 86.420 -31.940 86.870 -31.750 ;
        RECT 83.560 -32.170 86.870 -31.940 ;
        RECT 83.560 -32.250 84.020 -32.170 ;
        RECT 86.420 -32.260 86.870 -32.170 ;
        RECT 90.260 -31.520 90.710 -31.430 ;
        RECT 93.110 -31.520 93.570 -31.440 ;
        RECT 90.260 -31.750 93.570 -31.520 ;
        RECT 90.260 -31.940 90.710 -31.750 ;
        RECT 93.110 -31.940 93.570 -31.750 ;
        RECT 90.260 -32.170 93.570 -31.940 ;
        RECT 90.260 -32.260 90.710 -32.170 ;
        RECT 93.110 -32.250 93.570 -32.170 ;
        RECT 97.060 -31.520 97.520 -31.440 ;
        RECT 99.920 -31.520 100.370 -31.430 ;
        RECT 97.060 -31.750 100.370 -31.520 ;
        RECT 97.060 -31.940 97.520 -31.750 ;
        RECT 99.920 -31.940 100.370 -31.750 ;
        RECT 97.060 -32.170 100.370 -31.940 ;
        RECT 97.060 -32.250 97.520 -32.170 ;
        RECT 99.920 -32.260 100.370 -32.170 ;
        RECT 103.760 -31.520 104.210 -31.430 ;
        RECT 106.610 -31.520 107.070 -31.440 ;
        RECT 103.760 -31.750 107.070 -31.520 ;
        RECT 103.760 -31.940 104.210 -31.750 ;
        RECT 106.610 -31.940 107.070 -31.750 ;
        RECT 103.760 -32.170 107.070 -31.940 ;
        RECT 103.760 -32.260 104.210 -32.170 ;
        RECT 106.610 -32.250 107.070 -32.170 ;
        RECT 110.560 -31.520 111.020 -31.440 ;
        RECT 113.420 -31.520 113.870 -31.430 ;
        RECT 110.560 -31.750 113.870 -31.520 ;
        RECT 110.560 -31.940 111.020 -31.750 ;
        RECT 113.420 -31.940 113.870 -31.750 ;
        RECT 110.560 -32.170 113.870 -31.940 ;
        RECT 110.560 -32.250 111.020 -32.170 ;
        RECT 113.420 -32.260 113.870 -32.170 ;
        RECT 117.260 -31.520 117.710 -31.430 ;
        RECT 120.110 -31.520 120.570 -31.440 ;
        RECT 117.260 -31.750 120.570 -31.520 ;
        RECT 117.260 -31.940 117.710 -31.750 ;
        RECT 120.110 -31.940 120.570 -31.750 ;
        RECT 117.260 -32.170 120.570 -31.940 ;
        RECT 117.260 -32.260 117.710 -32.170 ;
        RECT 120.110 -32.250 120.570 -32.170 ;
        RECT 124.060 -31.520 124.520 -31.440 ;
        RECT 126.920 -31.520 127.370 -31.430 ;
        RECT 124.060 -31.750 127.370 -31.520 ;
        RECT 124.060 -31.940 124.520 -31.750 ;
        RECT 126.920 -31.940 127.370 -31.750 ;
        RECT 124.060 -32.170 127.370 -31.940 ;
        RECT 124.060 -32.250 124.520 -32.170 ;
        RECT 126.920 -32.260 127.370 -32.170 ;
        RECT 130.760 -31.520 131.210 -31.430 ;
        RECT 133.610 -31.520 134.070 -31.440 ;
        RECT 130.760 -31.750 134.070 -31.520 ;
        RECT 130.760 -31.940 131.210 -31.750 ;
        RECT 133.610 -31.940 134.070 -31.750 ;
        RECT 130.760 -32.170 134.070 -31.940 ;
        RECT 130.760 -32.260 131.210 -32.170 ;
        RECT 133.610 -32.250 134.070 -32.170 ;
        RECT 137.560 -31.520 138.020 -31.440 ;
        RECT 140.420 -31.520 140.870 -31.430 ;
        RECT 137.560 -31.750 140.870 -31.520 ;
        RECT 137.560 -31.940 138.020 -31.750 ;
        RECT 140.420 -31.940 140.870 -31.750 ;
        RECT 137.560 -32.170 140.870 -31.940 ;
        RECT 137.560 -32.250 138.020 -32.170 ;
        RECT 140.420 -32.260 140.870 -32.170 ;
        RECT 144.260 -31.520 144.710 -31.430 ;
        RECT 147.110 -31.520 147.570 -31.440 ;
        RECT 144.260 -31.750 147.570 -31.520 ;
        RECT 144.260 -31.940 144.710 -31.750 ;
        RECT 147.110 -31.940 147.570 -31.750 ;
        RECT 144.260 -32.170 147.570 -31.940 ;
        RECT 144.260 -32.260 144.710 -32.170 ;
        RECT 147.110 -32.250 147.570 -32.170 ;
        RECT 151.060 -31.520 151.520 -31.440 ;
        RECT 153.920 -31.520 154.370 -31.430 ;
        RECT 151.060 -31.750 154.370 -31.520 ;
        RECT 151.060 -31.940 151.520 -31.750 ;
        RECT 153.920 -31.940 154.370 -31.750 ;
        RECT 151.060 -32.170 154.370 -31.940 ;
        RECT 151.060 -32.250 151.520 -32.170 ;
        RECT 153.920 -32.260 154.370 -32.170 ;
        RECT 157.760 -31.520 158.210 -31.430 ;
        RECT 160.610 -31.520 161.070 -31.440 ;
        RECT 157.760 -31.750 161.070 -31.520 ;
        RECT 157.760 -31.940 158.210 -31.750 ;
        RECT 160.610 -31.940 161.070 -31.750 ;
        RECT 157.760 -32.170 161.070 -31.940 ;
        RECT 157.760 -32.260 158.210 -32.170 ;
        RECT 160.610 -32.250 161.070 -32.170 ;
        RECT 164.560 -31.520 165.020 -31.440 ;
        RECT 167.420 -31.520 167.870 -31.430 ;
        RECT 164.560 -31.750 167.870 -31.520 ;
        RECT 164.560 -31.940 165.020 -31.750 ;
        RECT 167.420 -31.940 167.870 -31.750 ;
        RECT 164.560 -32.170 167.870 -31.940 ;
        RECT 164.560 -32.250 165.020 -32.170 ;
        RECT 167.420 -32.260 167.870 -32.170 ;
        RECT 171.260 -31.520 171.710 -31.430 ;
        RECT 174.110 -31.520 174.570 -31.440 ;
        RECT 171.260 -31.750 174.570 -31.520 ;
        RECT 171.260 -31.940 171.710 -31.750 ;
        RECT 174.110 -31.940 174.570 -31.750 ;
        RECT 171.260 -32.170 174.570 -31.940 ;
        RECT 171.260 -32.260 171.710 -32.170 ;
        RECT 174.110 -32.250 174.570 -32.170 ;
        RECT 178.060 -31.520 178.520 -31.440 ;
        RECT 180.920 -31.520 181.370 -31.430 ;
        RECT 178.060 -31.750 181.370 -31.520 ;
        RECT 178.060 -31.940 178.520 -31.750 ;
        RECT 180.920 -31.940 181.370 -31.750 ;
        RECT 178.060 -32.170 181.370 -31.940 ;
        RECT 178.060 -32.250 178.520 -32.170 ;
        RECT 180.920 -32.260 181.370 -32.170 ;
        RECT 184.760 -31.520 185.210 -31.430 ;
        RECT 187.610 -31.520 188.070 -31.440 ;
        RECT 184.760 -31.750 188.070 -31.520 ;
        RECT 184.760 -31.940 185.210 -31.750 ;
        RECT 187.610 -31.940 188.070 -31.750 ;
        RECT 184.760 -32.170 188.070 -31.940 ;
        RECT 184.760 -32.260 185.210 -32.170 ;
        RECT 187.610 -32.250 188.070 -32.170 ;
        RECT 191.560 -31.520 192.020 -31.440 ;
        RECT 194.420 -31.520 194.870 -31.430 ;
        RECT 191.560 -31.750 194.870 -31.520 ;
        RECT 191.560 -31.940 192.020 -31.750 ;
        RECT 194.420 -31.940 194.870 -31.750 ;
        RECT 191.560 -32.170 194.870 -31.940 ;
        RECT 191.560 -32.250 192.020 -32.170 ;
        RECT 194.420 -32.260 194.870 -32.170 ;
        RECT 198.260 -31.520 198.710 -31.430 ;
        RECT 201.110 -31.520 201.570 -31.440 ;
        RECT 198.260 -31.750 201.570 -31.520 ;
        RECT 198.260 -31.940 198.710 -31.750 ;
        RECT 201.110 -31.940 201.570 -31.750 ;
        RECT 198.260 -32.170 201.570 -31.940 ;
        RECT 198.260 -32.260 198.710 -32.170 ;
        RECT 201.110 -32.250 201.570 -32.170 ;
        RECT 205.060 -31.520 205.520 -31.440 ;
        RECT 207.920 -31.520 208.370 -31.430 ;
        RECT 205.060 -31.750 208.370 -31.520 ;
        RECT 205.060 -31.940 205.520 -31.750 ;
        RECT 207.920 -31.940 208.370 -31.750 ;
        RECT 205.060 -32.170 208.370 -31.940 ;
        RECT 205.060 -32.250 205.520 -32.170 ;
        RECT 207.920 -32.260 208.370 -32.170 ;
        RECT 211.760 -31.520 212.210 -31.430 ;
        RECT 214.610 -31.520 215.070 -31.440 ;
        RECT 211.760 -31.750 215.070 -31.520 ;
        RECT 211.760 -31.940 212.210 -31.750 ;
        RECT 214.610 -31.940 215.070 -31.750 ;
        RECT 211.760 -32.170 215.070 -31.940 ;
        RECT 211.760 -32.260 212.210 -32.170 ;
        RECT 214.610 -32.250 215.070 -32.170 ;
        RECT 9.260 -35.130 9.710 -35.040 ;
        RECT 12.110 -35.130 12.570 -35.050 ;
        RECT 9.260 -35.360 12.570 -35.130 ;
        RECT 9.260 -35.550 9.710 -35.360 ;
        RECT 12.110 -35.550 12.570 -35.360 ;
        RECT 9.260 -35.780 12.570 -35.550 ;
        RECT 9.260 -35.870 9.710 -35.780 ;
        RECT 12.110 -35.860 12.570 -35.780 ;
        RECT 16.060 -35.130 16.520 -35.050 ;
        RECT 18.920 -35.130 19.370 -35.040 ;
        RECT 16.060 -35.360 19.370 -35.130 ;
        RECT 16.060 -35.550 16.520 -35.360 ;
        RECT 18.920 -35.550 19.370 -35.360 ;
        RECT 16.060 -35.780 19.370 -35.550 ;
        RECT 16.060 -35.860 16.520 -35.780 ;
        RECT 18.920 -35.870 19.370 -35.780 ;
        RECT 22.760 -35.130 23.210 -35.040 ;
        RECT 25.610 -35.130 26.070 -35.050 ;
        RECT 22.760 -35.360 26.070 -35.130 ;
        RECT 22.760 -35.550 23.210 -35.360 ;
        RECT 25.610 -35.550 26.070 -35.360 ;
        RECT 22.760 -35.780 26.070 -35.550 ;
        RECT 22.760 -35.870 23.210 -35.780 ;
        RECT 25.610 -35.860 26.070 -35.780 ;
        RECT 29.560 -35.130 30.020 -35.050 ;
        RECT 32.420 -35.130 32.870 -35.040 ;
        RECT 29.560 -35.360 32.870 -35.130 ;
        RECT 29.560 -35.550 30.020 -35.360 ;
        RECT 32.420 -35.550 32.870 -35.360 ;
        RECT 29.560 -35.780 32.870 -35.550 ;
        RECT 29.560 -35.860 30.020 -35.780 ;
        RECT 32.420 -35.870 32.870 -35.780 ;
        RECT 36.260 -35.130 36.710 -35.040 ;
        RECT 39.110 -35.130 39.570 -35.050 ;
        RECT 36.260 -35.360 39.570 -35.130 ;
        RECT 36.260 -35.550 36.710 -35.360 ;
        RECT 39.110 -35.550 39.570 -35.360 ;
        RECT 36.260 -35.780 39.570 -35.550 ;
        RECT 36.260 -35.870 36.710 -35.780 ;
        RECT 39.110 -35.860 39.570 -35.780 ;
        RECT 43.060 -35.130 43.520 -35.050 ;
        RECT 45.920 -35.130 46.370 -35.040 ;
        RECT 43.060 -35.360 46.370 -35.130 ;
        RECT 43.060 -35.550 43.520 -35.360 ;
        RECT 45.920 -35.550 46.370 -35.360 ;
        RECT 43.060 -35.780 46.370 -35.550 ;
        RECT 43.060 -35.860 43.520 -35.780 ;
        RECT 45.920 -35.870 46.370 -35.780 ;
        RECT 49.760 -35.130 50.210 -35.040 ;
        RECT 52.610 -35.130 53.070 -35.050 ;
        RECT 49.760 -35.360 53.070 -35.130 ;
        RECT 49.760 -35.550 50.210 -35.360 ;
        RECT 52.610 -35.550 53.070 -35.360 ;
        RECT 49.760 -35.780 53.070 -35.550 ;
        RECT 49.760 -35.870 50.210 -35.780 ;
        RECT 52.610 -35.860 53.070 -35.780 ;
        RECT 56.560 -35.130 57.020 -35.050 ;
        RECT 59.420 -35.130 59.870 -35.040 ;
        RECT 56.560 -35.360 59.870 -35.130 ;
        RECT 56.560 -35.550 57.020 -35.360 ;
        RECT 59.420 -35.550 59.870 -35.360 ;
        RECT 56.560 -35.780 59.870 -35.550 ;
        RECT 56.560 -35.860 57.020 -35.780 ;
        RECT 59.420 -35.870 59.870 -35.780 ;
        RECT 63.260 -35.130 63.710 -35.040 ;
        RECT 66.110 -35.130 66.570 -35.050 ;
        RECT 63.260 -35.360 66.570 -35.130 ;
        RECT 63.260 -35.550 63.710 -35.360 ;
        RECT 66.110 -35.550 66.570 -35.360 ;
        RECT 63.260 -35.780 66.570 -35.550 ;
        RECT 63.260 -35.870 63.710 -35.780 ;
        RECT 66.110 -35.860 66.570 -35.780 ;
        RECT 70.060 -35.130 70.520 -35.050 ;
        RECT 72.920 -35.130 73.370 -35.040 ;
        RECT 70.060 -35.360 73.370 -35.130 ;
        RECT 70.060 -35.550 70.520 -35.360 ;
        RECT 72.920 -35.550 73.370 -35.360 ;
        RECT 70.060 -35.780 73.370 -35.550 ;
        RECT 70.060 -35.860 70.520 -35.780 ;
        RECT 72.920 -35.870 73.370 -35.780 ;
        RECT 76.760 -35.130 77.210 -35.040 ;
        RECT 79.610 -35.130 80.070 -35.050 ;
        RECT 76.760 -35.360 80.070 -35.130 ;
        RECT 76.760 -35.550 77.210 -35.360 ;
        RECT 79.610 -35.550 80.070 -35.360 ;
        RECT 76.760 -35.780 80.070 -35.550 ;
        RECT 76.760 -35.870 77.210 -35.780 ;
        RECT 79.610 -35.860 80.070 -35.780 ;
        RECT 83.560 -35.130 84.020 -35.050 ;
        RECT 86.420 -35.130 86.870 -35.040 ;
        RECT 83.560 -35.360 86.870 -35.130 ;
        RECT 83.560 -35.550 84.020 -35.360 ;
        RECT 86.420 -35.550 86.870 -35.360 ;
        RECT 83.560 -35.780 86.870 -35.550 ;
        RECT 83.560 -35.860 84.020 -35.780 ;
        RECT 86.420 -35.870 86.870 -35.780 ;
        RECT 90.260 -35.130 90.710 -35.040 ;
        RECT 93.110 -35.130 93.570 -35.050 ;
        RECT 90.260 -35.360 93.570 -35.130 ;
        RECT 90.260 -35.550 90.710 -35.360 ;
        RECT 93.110 -35.550 93.570 -35.360 ;
        RECT 90.260 -35.780 93.570 -35.550 ;
        RECT 90.260 -35.870 90.710 -35.780 ;
        RECT 93.110 -35.860 93.570 -35.780 ;
        RECT 97.060 -35.130 97.520 -35.050 ;
        RECT 99.920 -35.130 100.370 -35.040 ;
        RECT 97.060 -35.360 100.370 -35.130 ;
        RECT 97.060 -35.550 97.520 -35.360 ;
        RECT 99.920 -35.550 100.370 -35.360 ;
        RECT 97.060 -35.780 100.370 -35.550 ;
        RECT 97.060 -35.860 97.520 -35.780 ;
        RECT 99.920 -35.870 100.370 -35.780 ;
        RECT 103.760 -35.130 104.210 -35.040 ;
        RECT 106.610 -35.130 107.070 -35.050 ;
        RECT 103.760 -35.360 107.070 -35.130 ;
        RECT 103.760 -35.550 104.210 -35.360 ;
        RECT 106.610 -35.550 107.070 -35.360 ;
        RECT 103.760 -35.780 107.070 -35.550 ;
        RECT 103.760 -35.870 104.210 -35.780 ;
        RECT 106.610 -35.860 107.070 -35.780 ;
        RECT 110.560 -35.130 111.020 -35.050 ;
        RECT 113.420 -35.130 113.870 -35.040 ;
        RECT 110.560 -35.360 113.870 -35.130 ;
        RECT 110.560 -35.550 111.020 -35.360 ;
        RECT 113.420 -35.550 113.870 -35.360 ;
        RECT 110.560 -35.780 113.870 -35.550 ;
        RECT 110.560 -35.860 111.020 -35.780 ;
        RECT 113.420 -35.870 113.870 -35.780 ;
        RECT 117.260 -35.130 117.710 -35.040 ;
        RECT 120.110 -35.130 120.570 -35.050 ;
        RECT 117.260 -35.360 120.570 -35.130 ;
        RECT 117.260 -35.550 117.710 -35.360 ;
        RECT 120.110 -35.550 120.570 -35.360 ;
        RECT 117.260 -35.780 120.570 -35.550 ;
        RECT 117.260 -35.870 117.710 -35.780 ;
        RECT 120.110 -35.860 120.570 -35.780 ;
        RECT 124.060 -35.130 124.520 -35.050 ;
        RECT 126.920 -35.130 127.370 -35.040 ;
        RECT 124.060 -35.360 127.370 -35.130 ;
        RECT 124.060 -35.550 124.520 -35.360 ;
        RECT 126.920 -35.550 127.370 -35.360 ;
        RECT 124.060 -35.780 127.370 -35.550 ;
        RECT 124.060 -35.860 124.520 -35.780 ;
        RECT 126.920 -35.870 127.370 -35.780 ;
        RECT 130.760 -35.130 131.210 -35.040 ;
        RECT 133.610 -35.130 134.070 -35.050 ;
        RECT 130.760 -35.360 134.070 -35.130 ;
        RECT 130.760 -35.550 131.210 -35.360 ;
        RECT 133.610 -35.550 134.070 -35.360 ;
        RECT 130.760 -35.780 134.070 -35.550 ;
        RECT 130.760 -35.870 131.210 -35.780 ;
        RECT 133.610 -35.860 134.070 -35.780 ;
        RECT 137.560 -35.130 138.020 -35.050 ;
        RECT 140.420 -35.130 140.870 -35.040 ;
        RECT 137.560 -35.360 140.870 -35.130 ;
        RECT 137.560 -35.550 138.020 -35.360 ;
        RECT 140.420 -35.550 140.870 -35.360 ;
        RECT 137.560 -35.780 140.870 -35.550 ;
        RECT 137.560 -35.860 138.020 -35.780 ;
        RECT 140.420 -35.870 140.870 -35.780 ;
        RECT 144.260 -35.130 144.710 -35.040 ;
        RECT 147.110 -35.130 147.570 -35.050 ;
        RECT 144.260 -35.360 147.570 -35.130 ;
        RECT 144.260 -35.550 144.710 -35.360 ;
        RECT 147.110 -35.550 147.570 -35.360 ;
        RECT 144.260 -35.780 147.570 -35.550 ;
        RECT 144.260 -35.870 144.710 -35.780 ;
        RECT 147.110 -35.860 147.570 -35.780 ;
        RECT 151.060 -35.130 151.520 -35.050 ;
        RECT 153.920 -35.130 154.370 -35.040 ;
        RECT 151.060 -35.360 154.370 -35.130 ;
        RECT 151.060 -35.550 151.520 -35.360 ;
        RECT 153.920 -35.550 154.370 -35.360 ;
        RECT 151.060 -35.780 154.370 -35.550 ;
        RECT 151.060 -35.860 151.520 -35.780 ;
        RECT 153.920 -35.870 154.370 -35.780 ;
        RECT 157.760 -35.130 158.210 -35.040 ;
        RECT 160.610 -35.130 161.070 -35.050 ;
        RECT 157.760 -35.360 161.070 -35.130 ;
        RECT 157.760 -35.550 158.210 -35.360 ;
        RECT 160.610 -35.550 161.070 -35.360 ;
        RECT 157.760 -35.780 161.070 -35.550 ;
        RECT 157.760 -35.870 158.210 -35.780 ;
        RECT 160.610 -35.860 161.070 -35.780 ;
        RECT 164.560 -35.130 165.020 -35.050 ;
        RECT 167.420 -35.130 167.870 -35.040 ;
        RECT 164.560 -35.360 167.870 -35.130 ;
        RECT 164.560 -35.550 165.020 -35.360 ;
        RECT 167.420 -35.550 167.870 -35.360 ;
        RECT 164.560 -35.780 167.870 -35.550 ;
        RECT 164.560 -35.860 165.020 -35.780 ;
        RECT 167.420 -35.870 167.870 -35.780 ;
        RECT 171.260 -35.130 171.710 -35.040 ;
        RECT 174.110 -35.130 174.570 -35.050 ;
        RECT 171.260 -35.360 174.570 -35.130 ;
        RECT 171.260 -35.550 171.710 -35.360 ;
        RECT 174.110 -35.550 174.570 -35.360 ;
        RECT 171.260 -35.780 174.570 -35.550 ;
        RECT 171.260 -35.870 171.710 -35.780 ;
        RECT 174.110 -35.860 174.570 -35.780 ;
        RECT 178.060 -35.130 178.520 -35.050 ;
        RECT 180.920 -35.130 181.370 -35.040 ;
        RECT 178.060 -35.360 181.370 -35.130 ;
        RECT 178.060 -35.550 178.520 -35.360 ;
        RECT 180.920 -35.550 181.370 -35.360 ;
        RECT 178.060 -35.780 181.370 -35.550 ;
        RECT 178.060 -35.860 178.520 -35.780 ;
        RECT 180.920 -35.870 181.370 -35.780 ;
        RECT 184.760 -35.130 185.210 -35.040 ;
        RECT 187.610 -35.130 188.070 -35.050 ;
        RECT 184.760 -35.360 188.070 -35.130 ;
        RECT 184.760 -35.550 185.210 -35.360 ;
        RECT 187.610 -35.550 188.070 -35.360 ;
        RECT 184.760 -35.780 188.070 -35.550 ;
        RECT 184.760 -35.870 185.210 -35.780 ;
        RECT 187.610 -35.860 188.070 -35.780 ;
        RECT 191.560 -35.130 192.020 -35.050 ;
        RECT 194.420 -35.130 194.870 -35.040 ;
        RECT 191.560 -35.360 194.870 -35.130 ;
        RECT 191.560 -35.550 192.020 -35.360 ;
        RECT 194.420 -35.550 194.870 -35.360 ;
        RECT 191.560 -35.780 194.870 -35.550 ;
        RECT 191.560 -35.860 192.020 -35.780 ;
        RECT 194.420 -35.870 194.870 -35.780 ;
        RECT 198.260 -35.130 198.710 -35.040 ;
        RECT 201.110 -35.130 201.570 -35.050 ;
        RECT 198.260 -35.360 201.570 -35.130 ;
        RECT 198.260 -35.550 198.710 -35.360 ;
        RECT 201.110 -35.550 201.570 -35.360 ;
        RECT 198.260 -35.780 201.570 -35.550 ;
        RECT 198.260 -35.870 198.710 -35.780 ;
        RECT 201.110 -35.860 201.570 -35.780 ;
        RECT 205.060 -35.130 205.520 -35.050 ;
        RECT 207.920 -35.130 208.370 -35.040 ;
        RECT 205.060 -35.360 208.370 -35.130 ;
        RECT 205.060 -35.550 205.520 -35.360 ;
        RECT 207.920 -35.550 208.370 -35.360 ;
        RECT 205.060 -35.780 208.370 -35.550 ;
        RECT 205.060 -35.860 205.520 -35.780 ;
        RECT 207.920 -35.870 208.370 -35.780 ;
        RECT 211.760 -35.130 212.210 -35.040 ;
        RECT 214.610 -35.130 215.070 -35.050 ;
        RECT 211.760 -35.360 215.070 -35.130 ;
        RECT 211.760 -35.550 212.210 -35.360 ;
        RECT 214.610 -35.550 215.070 -35.360 ;
        RECT 211.760 -35.780 215.070 -35.550 ;
        RECT 211.760 -35.870 212.210 -35.780 ;
        RECT 214.610 -35.860 215.070 -35.780 ;
        RECT 9.260 -38.740 9.710 -38.650 ;
        RECT 12.110 -38.740 12.570 -38.660 ;
        RECT 9.260 -38.970 12.570 -38.740 ;
        RECT 9.260 -39.160 9.710 -38.970 ;
        RECT 12.110 -39.160 12.570 -38.970 ;
        RECT 9.260 -39.390 12.570 -39.160 ;
        RECT 9.260 -39.480 9.710 -39.390 ;
        RECT 12.110 -39.470 12.570 -39.390 ;
        RECT 16.060 -38.740 16.520 -38.660 ;
        RECT 18.920 -38.740 19.370 -38.650 ;
        RECT 16.060 -38.970 19.370 -38.740 ;
        RECT 16.060 -39.160 16.520 -38.970 ;
        RECT 18.920 -39.160 19.370 -38.970 ;
        RECT 16.060 -39.390 19.370 -39.160 ;
        RECT 16.060 -39.470 16.520 -39.390 ;
        RECT 18.920 -39.480 19.370 -39.390 ;
        RECT 22.760 -38.740 23.210 -38.650 ;
        RECT 25.610 -38.740 26.070 -38.660 ;
        RECT 22.760 -38.970 26.070 -38.740 ;
        RECT 22.760 -39.160 23.210 -38.970 ;
        RECT 25.610 -39.160 26.070 -38.970 ;
        RECT 22.760 -39.390 26.070 -39.160 ;
        RECT 22.760 -39.480 23.210 -39.390 ;
        RECT 25.610 -39.470 26.070 -39.390 ;
        RECT 29.560 -38.740 30.020 -38.660 ;
        RECT 32.420 -38.740 32.870 -38.650 ;
        RECT 29.560 -38.970 32.870 -38.740 ;
        RECT 29.560 -39.160 30.020 -38.970 ;
        RECT 32.420 -39.160 32.870 -38.970 ;
        RECT 29.560 -39.390 32.870 -39.160 ;
        RECT 29.560 -39.470 30.020 -39.390 ;
        RECT 32.420 -39.480 32.870 -39.390 ;
        RECT 36.260 -38.740 36.710 -38.650 ;
        RECT 39.110 -38.740 39.570 -38.660 ;
        RECT 36.260 -38.970 39.570 -38.740 ;
        RECT 36.260 -39.160 36.710 -38.970 ;
        RECT 39.110 -39.160 39.570 -38.970 ;
        RECT 36.260 -39.390 39.570 -39.160 ;
        RECT 36.260 -39.480 36.710 -39.390 ;
        RECT 39.110 -39.470 39.570 -39.390 ;
        RECT 43.060 -38.740 43.520 -38.660 ;
        RECT 45.920 -38.740 46.370 -38.650 ;
        RECT 43.060 -38.970 46.370 -38.740 ;
        RECT 43.060 -39.160 43.520 -38.970 ;
        RECT 45.920 -39.160 46.370 -38.970 ;
        RECT 43.060 -39.390 46.370 -39.160 ;
        RECT 43.060 -39.470 43.520 -39.390 ;
        RECT 45.920 -39.480 46.370 -39.390 ;
        RECT 49.760 -38.740 50.210 -38.650 ;
        RECT 52.610 -38.740 53.070 -38.660 ;
        RECT 49.760 -38.970 53.070 -38.740 ;
        RECT 49.760 -39.160 50.210 -38.970 ;
        RECT 52.610 -39.160 53.070 -38.970 ;
        RECT 49.760 -39.390 53.070 -39.160 ;
        RECT 49.760 -39.480 50.210 -39.390 ;
        RECT 52.610 -39.470 53.070 -39.390 ;
        RECT 56.560 -38.740 57.020 -38.660 ;
        RECT 59.420 -38.740 59.870 -38.650 ;
        RECT 56.560 -38.970 59.870 -38.740 ;
        RECT 56.560 -39.160 57.020 -38.970 ;
        RECT 59.420 -39.160 59.870 -38.970 ;
        RECT 56.560 -39.390 59.870 -39.160 ;
        RECT 56.560 -39.470 57.020 -39.390 ;
        RECT 59.420 -39.480 59.870 -39.390 ;
        RECT 63.260 -38.740 63.710 -38.650 ;
        RECT 66.110 -38.740 66.570 -38.660 ;
        RECT 63.260 -38.970 66.570 -38.740 ;
        RECT 63.260 -39.160 63.710 -38.970 ;
        RECT 66.110 -39.160 66.570 -38.970 ;
        RECT 63.260 -39.390 66.570 -39.160 ;
        RECT 63.260 -39.480 63.710 -39.390 ;
        RECT 66.110 -39.470 66.570 -39.390 ;
        RECT 70.060 -38.740 70.520 -38.660 ;
        RECT 72.920 -38.740 73.370 -38.650 ;
        RECT 70.060 -38.970 73.370 -38.740 ;
        RECT 70.060 -39.160 70.520 -38.970 ;
        RECT 72.920 -39.160 73.370 -38.970 ;
        RECT 70.060 -39.390 73.370 -39.160 ;
        RECT 70.060 -39.470 70.520 -39.390 ;
        RECT 72.920 -39.480 73.370 -39.390 ;
        RECT 76.760 -38.740 77.210 -38.650 ;
        RECT 79.610 -38.740 80.070 -38.660 ;
        RECT 76.760 -38.970 80.070 -38.740 ;
        RECT 76.760 -39.160 77.210 -38.970 ;
        RECT 79.610 -39.160 80.070 -38.970 ;
        RECT 76.760 -39.390 80.070 -39.160 ;
        RECT 76.760 -39.480 77.210 -39.390 ;
        RECT 79.610 -39.470 80.070 -39.390 ;
        RECT 83.560 -38.740 84.020 -38.660 ;
        RECT 86.420 -38.740 86.870 -38.650 ;
        RECT 83.560 -38.970 86.870 -38.740 ;
        RECT 83.560 -39.160 84.020 -38.970 ;
        RECT 86.420 -39.160 86.870 -38.970 ;
        RECT 83.560 -39.390 86.870 -39.160 ;
        RECT 83.560 -39.470 84.020 -39.390 ;
        RECT 86.420 -39.480 86.870 -39.390 ;
        RECT 90.260 -38.740 90.710 -38.650 ;
        RECT 93.110 -38.740 93.570 -38.660 ;
        RECT 90.260 -38.970 93.570 -38.740 ;
        RECT 90.260 -39.160 90.710 -38.970 ;
        RECT 93.110 -39.160 93.570 -38.970 ;
        RECT 90.260 -39.390 93.570 -39.160 ;
        RECT 90.260 -39.480 90.710 -39.390 ;
        RECT 93.110 -39.470 93.570 -39.390 ;
        RECT 97.060 -38.740 97.520 -38.660 ;
        RECT 99.920 -38.740 100.370 -38.650 ;
        RECT 97.060 -38.970 100.370 -38.740 ;
        RECT 97.060 -39.160 97.520 -38.970 ;
        RECT 99.920 -39.160 100.370 -38.970 ;
        RECT 97.060 -39.390 100.370 -39.160 ;
        RECT 97.060 -39.470 97.520 -39.390 ;
        RECT 99.920 -39.480 100.370 -39.390 ;
        RECT 103.760 -38.740 104.210 -38.650 ;
        RECT 106.610 -38.740 107.070 -38.660 ;
        RECT 103.760 -38.970 107.070 -38.740 ;
        RECT 103.760 -39.160 104.210 -38.970 ;
        RECT 106.610 -39.160 107.070 -38.970 ;
        RECT 103.760 -39.390 107.070 -39.160 ;
        RECT 103.760 -39.480 104.210 -39.390 ;
        RECT 106.610 -39.470 107.070 -39.390 ;
        RECT 110.560 -38.740 111.020 -38.660 ;
        RECT 113.420 -38.740 113.870 -38.650 ;
        RECT 110.560 -38.970 113.870 -38.740 ;
        RECT 110.560 -39.160 111.020 -38.970 ;
        RECT 113.420 -39.160 113.870 -38.970 ;
        RECT 110.560 -39.390 113.870 -39.160 ;
        RECT 110.560 -39.470 111.020 -39.390 ;
        RECT 113.420 -39.480 113.870 -39.390 ;
        RECT 117.260 -38.740 117.710 -38.650 ;
        RECT 120.110 -38.740 120.570 -38.660 ;
        RECT 117.260 -38.970 120.570 -38.740 ;
        RECT 117.260 -39.160 117.710 -38.970 ;
        RECT 120.110 -39.160 120.570 -38.970 ;
        RECT 117.260 -39.390 120.570 -39.160 ;
        RECT 117.260 -39.480 117.710 -39.390 ;
        RECT 120.110 -39.470 120.570 -39.390 ;
        RECT 124.060 -38.740 124.520 -38.660 ;
        RECT 126.920 -38.740 127.370 -38.650 ;
        RECT 124.060 -38.970 127.370 -38.740 ;
        RECT 124.060 -39.160 124.520 -38.970 ;
        RECT 126.920 -39.160 127.370 -38.970 ;
        RECT 124.060 -39.390 127.370 -39.160 ;
        RECT 124.060 -39.470 124.520 -39.390 ;
        RECT 126.920 -39.480 127.370 -39.390 ;
        RECT 130.760 -38.740 131.210 -38.650 ;
        RECT 133.610 -38.740 134.070 -38.660 ;
        RECT 130.760 -38.970 134.070 -38.740 ;
        RECT 130.760 -39.160 131.210 -38.970 ;
        RECT 133.610 -39.160 134.070 -38.970 ;
        RECT 130.760 -39.390 134.070 -39.160 ;
        RECT 130.760 -39.480 131.210 -39.390 ;
        RECT 133.610 -39.470 134.070 -39.390 ;
        RECT 137.560 -38.740 138.020 -38.660 ;
        RECT 140.420 -38.740 140.870 -38.650 ;
        RECT 137.560 -38.970 140.870 -38.740 ;
        RECT 137.560 -39.160 138.020 -38.970 ;
        RECT 140.420 -39.160 140.870 -38.970 ;
        RECT 137.560 -39.390 140.870 -39.160 ;
        RECT 137.560 -39.470 138.020 -39.390 ;
        RECT 140.420 -39.480 140.870 -39.390 ;
        RECT 144.260 -38.740 144.710 -38.650 ;
        RECT 147.110 -38.740 147.570 -38.660 ;
        RECT 144.260 -38.970 147.570 -38.740 ;
        RECT 144.260 -39.160 144.710 -38.970 ;
        RECT 147.110 -39.160 147.570 -38.970 ;
        RECT 144.260 -39.390 147.570 -39.160 ;
        RECT 144.260 -39.480 144.710 -39.390 ;
        RECT 147.110 -39.470 147.570 -39.390 ;
        RECT 151.060 -38.740 151.520 -38.660 ;
        RECT 153.920 -38.740 154.370 -38.650 ;
        RECT 151.060 -38.970 154.370 -38.740 ;
        RECT 151.060 -39.160 151.520 -38.970 ;
        RECT 153.920 -39.160 154.370 -38.970 ;
        RECT 151.060 -39.390 154.370 -39.160 ;
        RECT 151.060 -39.470 151.520 -39.390 ;
        RECT 153.920 -39.480 154.370 -39.390 ;
        RECT 157.760 -38.740 158.210 -38.650 ;
        RECT 160.610 -38.740 161.070 -38.660 ;
        RECT 157.760 -38.970 161.070 -38.740 ;
        RECT 157.760 -39.160 158.210 -38.970 ;
        RECT 160.610 -39.160 161.070 -38.970 ;
        RECT 157.760 -39.390 161.070 -39.160 ;
        RECT 157.760 -39.480 158.210 -39.390 ;
        RECT 160.610 -39.470 161.070 -39.390 ;
        RECT 164.560 -38.740 165.020 -38.660 ;
        RECT 167.420 -38.740 167.870 -38.650 ;
        RECT 164.560 -38.970 167.870 -38.740 ;
        RECT 164.560 -39.160 165.020 -38.970 ;
        RECT 167.420 -39.160 167.870 -38.970 ;
        RECT 164.560 -39.390 167.870 -39.160 ;
        RECT 164.560 -39.470 165.020 -39.390 ;
        RECT 167.420 -39.480 167.870 -39.390 ;
        RECT 171.260 -38.740 171.710 -38.650 ;
        RECT 174.110 -38.740 174.570 -38.660 ;
        RECT 171.260 -38.970 174.570 -38.740 ;
        RECT 171.260 -39.160 171.710 -38.970 ;
        RECT 174.110 -39.160 174.570 -38.970 ;
        RECT 171.260 -39.390 174.570 -39.160 ;
        RECT 171.260 -39.480 171.710 -39.390 ;
        RECT 174.110 -39.470 174.570 -39.390 ;
        RECT 178.060 -38.740 178.520 -38.660 ;
        RECT 180.920 -38.740 181.370 -38.650 ;
        RECT 178.060 -38.970 181.370 -38.740 ;
        RECT 178.060 -39.160 178.520 -38.970 ;
        RECT 180.920 -39.160 181.370 -38.970 ;
        RECT 178.060 -39.390 181.370 -39.160 ;
        RECT 178.060 -39.470 178.520 -39.390 ;
        RECT 180.920 -39.480 181.370 -39.390 ;
        RECT 184.760 -38.740 185.210 -38.650 ;
        RECT 187.610 -38.740 188.070 -38.660 ;
        RECT 184.760 -38.970 188.070 -38.740 ;
        RECT 184.760 -39.160 185.210 -38.970 ;
        RECT 187.610 -39.160 188.070 -38.970 ;
        RECT 184.760 -39.390 188.070 -39.160 ;
        RECT 184.760 -39.480 185.210 -39.390 ;
        RECT 187.610 -39.470 188.070 -39.390 ;
        RECT 191.560 -38.740 192.020 -38.660 ;
        RECT 194.420 -38.740 194.870 -38.650 ;
        RECT 191.560 -38.970 194.870 -38.740 ;
        RECT 191.560 -39.160 192.020 -38.970 ;
        RECT 194.420 -39.160 194.870 -38.970 ;
        RECT 191.560 -39.390 194.870 -39.160 ;
        RECT 191.560 -39.470 192.020 -39.390 ;
        RECT 194.420 -39.480 194.870 -39.390 ;
        RECT 198.260 -38.740 198.710 -38.650 ;
        RECT 201.110 -38.740 201.570 -38.660 ;
        RECT 198.260 -38.970 201.570 -38.740 ;
        RECT 198.260 -39.160 198.710 -38.970 ;
        RECT 201.110 -39.160 201.570 -38.970 ;
        RECT 198.260 -39.390 201.570 -39.160 ;
        RECT 198.260 -39.480 198.710 -39.390 ;
        RECT 201.110 -39.470 201.570 -39.390 ;
        RECT 205.060 -38.740 205.520 -38.660 ;
        RECT 207.920 -38.740 208.370 -38.650 ;
        RECT 205.060 -38.970 208.370 -38.740 ;
        RECT 205.060 -39.160 205.520 -38.970 ;
        RECT 207.920 -39.160 208.370 -38.970 ;
        RECT 205.060 -39.390 208.370 -39.160 ;
        RECT 205.060 -39.470 205.520 -39.390 ;
        RECT 207.920 -39.480 208.370 -39.390 ;
        RECT 211.760 -38.740 212.210 -38.650 ;
        RECT 214.610 -38.740 215.070 -38.660 ;
        RECT 211.760 -38.970 215.070 -38.740 ;
        RECT 211.760 -39.160 212.210 -38.970 ;
        RECT 214.610 -39.160 215.070 -38.970 ;
        RECT 211.760 -39.390 215.070 -39.160 ;
        RECT 211.760 -39.480 212.210 -39.390 ;
        RECT 214.610 -39.470 215.070 -39.390 ;
  END
END IMPACTSram
END LIBRARY

