// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0


module BankWordDecoder (
`ifdef USE_POWER_PINS
    inout vccd1,	// User area 1 1.8V supply
    inout vssd1,	// User area 1 digital ground
`endif
	input clk,
	input [9:0] sel,
	output reg [1023:0] address

);

    integer i;
    always@(posedge clk) begin
	 address[0] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[1] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[2] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[3] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[4] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[5] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[6] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[7] = sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[8] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[9] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[10] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[11] = sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[12] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[13] = sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[14] = ~sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[15] = sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[16] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[17] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[18] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[19] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[20] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[21] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[22] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[23] = sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[24] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[25] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[26] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[27] = sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[28] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[29] = sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[30] = ~sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[31] = sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[32] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[33] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[34] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[35] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[36] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[37] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[38] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[39] = sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[40] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[41] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[42] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[43] = sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[44] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[45] = sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[46] = ~sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[47] = sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[48] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[49] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[50] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[51] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[52] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[53] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[54] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[55] = sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[56] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[57] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[58] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[59] = sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[60] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[61] = sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[62] = ~sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[63] = sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[64] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[65] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[66] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[67] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[68] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[69] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[70] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[71] = sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[72] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[73] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[74] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[75] = sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[76] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[77] = sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[78] = ~sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[79] = sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[80] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[81] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[82] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[83] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[84] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[85] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[86] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[87] = sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[88] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[89] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[90] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[91] = sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[92] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[93] = sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[94] = ~sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[95] = sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[96] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[97] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[98] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[99] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[100] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[101] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[102] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[103] = sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[104] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[105] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[106] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[107] = sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[108] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[109] = sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[110] = ~sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[111] = sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[112] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[113] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[114] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[115] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[116] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[117] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[118] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[119] = sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[120] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[121] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[122] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[123] = sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[124] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[125] = sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[126] = ~sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[127] = sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
	 address[128] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[129] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[130] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[131] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[132] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[133] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[134] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[135] = sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[136] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[137] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[138] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[139] = sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[140] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[141] = sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[142] = ~sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[143] = sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[144] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[145] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[146] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[147] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[148] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[149] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[150] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[151] = sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[152] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[153] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[154] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[155] = sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[156] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[157] = sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[158] = ~sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[159] = sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[160] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[161] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[162] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[163] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[164] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[165] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[166] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[167] = sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[168] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[169] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[170] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[171] = sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[172] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[173] = sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[174] = ~sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[175] = sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[176] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[177] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[178] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[179] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[180] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[181] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[182] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[183] = sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[184] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[185] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[186] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[187] = sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[188] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[189] = sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[190] = ~sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[191] = sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[192] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[193] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[194] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[195] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[196] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[197] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[198] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[199] = sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[200] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[201] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[202] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[203] = sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[204] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[205] = sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[206] = ~sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[207] = sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[208] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[209] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[210] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[211] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[212] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[213] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[214] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[215] = sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[216] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[217] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[218] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[219] = sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[220] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[221] = sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[222] = ~sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[223] = sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[224] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[225] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[226] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[227] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[228] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[229] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[230] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[231] = sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[232] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[233] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[234] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[235] = sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[236] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[237] = sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[238] = ~sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[239] = sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[240] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[241] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[242] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[243] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[244] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[245] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[246] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[247] = sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[248] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[249] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[250] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[251] = sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[252] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[253] = sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[254] = ~sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[255] = sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
	 address[256] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[257] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[258] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[259] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[260] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[261] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[262] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[263] = sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[264] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[265] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[266] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[267] = sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[268] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[269] = sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[270] = ~sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[271] = sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[272] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[273] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[274] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[275] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[276] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[277] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[278] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[279] = sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[280] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[281] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[282] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[283] = sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[284] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[285] = sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[286] = ~sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[287] = sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[288] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[289] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[290] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[291] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[292] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[293] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[294] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[295] = sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[296] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[297] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[298] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[299] = sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[300] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[301] = sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[302] = ~sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[303] = sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[304] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[305] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[306] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[307] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[308] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[309] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[310] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[311] = sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[312] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[313] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[314] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[315] = sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[316] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[317] = sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[318] = ~sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[319] = sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[320] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[321] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[322] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[323] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[324] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[325] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[326] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[327] = sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[328] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[329] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[330] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[331] = sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[332] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[333] = sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[334] = ~sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[335] = sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[336] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[337] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[338] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[339] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[340] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[341] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[342] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[343] = sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[344] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[345] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[346] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[347] = sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[348] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[349] = sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[350] = ~sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[351] = sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[352] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[353] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[354] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[355] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[356] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[357] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[358] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[359] = sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[360] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[361] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[362] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[363] = sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[364] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[365] = sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[366] = ~sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[367] = sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[368] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[369] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[370] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[371] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[372] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[373] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[374] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[375] = sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[376] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[377] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[378] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[379] = sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[380] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[381] = sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[382] = ~sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[383] = sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
	 address[384] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[385] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[386] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[387] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[388] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[389] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[390] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[391] = sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[392] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[393] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[394] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[395] = sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[396] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[397] = sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[398] = ~sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[399] = sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[400] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[401] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[402] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[403] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[404] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[405] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[406] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[407] = sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[408] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[409] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[410] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[411] = sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[412] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[413] = sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[414] = ~sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[415] = sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[416] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[417] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[418] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[419] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[420] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[421] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[422] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[423] = sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[424] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[425] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[426] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[427] = sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[428] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[429] = sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[430] = ~sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[431] = sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[432] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[433] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[434] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[435] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[436] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[437] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[438] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[439] = sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[440] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[441] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[442] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[443] = sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[444] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[445] = sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[446] = ~sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[447] = sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[448] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[449] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[450] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[451] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[452] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[453] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[454] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[455] = sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[456] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[457] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[458] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[459] = sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[460] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[461] = sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[462] = ~sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[463] = sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[464] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[465] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[466] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[467] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[468] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[469] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[470] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[471] = sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[472] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[473] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[474] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[475] = sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[476] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[477] = sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[478] = ~sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[479] = sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[480] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[481] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[482] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[483] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[484] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[485] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[486] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[487] = sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[488] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[489] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[490] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[491] = sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[492] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[493] = sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[494] = ~sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[495] = sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[496] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[497] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[498] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[499] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[500] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[501] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[502] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[503] = sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[504] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[505] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[506] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[507] = sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[508] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[509] = sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[510] = ~sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[511] = sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
	 address[512] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[513] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[514] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[515] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[516] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[517] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[518] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[519] = sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[520] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[521] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[522] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[523] = sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[524] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[525] = sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[526] = ~sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[527] = sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[528] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[529] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[530] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[531] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[532] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[533] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[534] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[535] = sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[536] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[537] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[538] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[539] = sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[540] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[541] = sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[542] = ~sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[543] = sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[544] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[545] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[546] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[547] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[548] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[549] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[550] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[551] = sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[552] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[553] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[554] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[555] = sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[556] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[557] = sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[558] = ~sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[559] = sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[560] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[561] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[562] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[563] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[564] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[565] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[566] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[567] = sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[568] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[569] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[570] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[571] = sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[572] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[573] = sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[574] = ~sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[575] = sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[576] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[577] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[578] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[579] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[580] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[581] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[582] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[583] = sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[584] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[585] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[586] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[587] = sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[588] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[589] = sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[590] = ~sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[591] = sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[592] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[593] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[594] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[595] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[596] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[597] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[598] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[599] = sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[600] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[601] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[602] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[603] = sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[604] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[605] = sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[606] = ~sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[607] = sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[608] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[609] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[610] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[611] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[612] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[613] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[614] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[615] = sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[616] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[617] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[618] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[619] = sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[620] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[621] = sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[622] = ~sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[623] = sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[624] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[625] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[626] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[627] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[628] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[629] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[630] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[631] = sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[632] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[633] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[634] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[635] = sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[636] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[637] = sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[638] = ~sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[639] = sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
	 address[640] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[641] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[642] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[643] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[644] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[645] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[646] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[647] = sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[648] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[649] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[650] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[651] = sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[652] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[653] = sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[654] = ~sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[655] = sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[656] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[657] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[658] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[659] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[660] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[661] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[662] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[663] = sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[664] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[665] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[666] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[667] = sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[668] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[669] = sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[670] = ~sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[671] = sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[672] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[673] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[674] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[675] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[676] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[677] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[678] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[679] = sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[680] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[681] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[682] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[683] = sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[684] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[685] = sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[686] = ~sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[687] = sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[688] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[689] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[690] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[691] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[692] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[693] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[694] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[695] = sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[696] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[697] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[698] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[699] = sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[700] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[701] = sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[702] = ~sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[703] = sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[704] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[705] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[706] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[707] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[708] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[709] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[710] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[711] = sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[712] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[713] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[714] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[715] = sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[716] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[717] = sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[718] = ~sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[719] = sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[720] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[721] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[722] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[723] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[724] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[725] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[726] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[727] = sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[728] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[729] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[730] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[731] = sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[732] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[733] = sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[734] = ~sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[735] = sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[736] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[737] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[738] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[739] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[740] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[741] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[742] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[743] = sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[744] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[745] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[746] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[747] = sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[748] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[749] = sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[750] = ~sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[751] = sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[752] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[753] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[754] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[755] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[756] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[757] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[758] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[759] = sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[760] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[761] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[762] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[763] = sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[764] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[765] = sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[766] = ~sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[767] = sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
	 address[768] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[769] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[770] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[771] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[772] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[773] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[774] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[775] = sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[776] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[777] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[778] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[779] = sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[780] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[781] = sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[782] = ~sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[783] = sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[784] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[785] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[786] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[787] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[788] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[789] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[790] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[791] = sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[792] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[793] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[794] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[795] = sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[796] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[797] = sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[798] = ~sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[799] = sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[800] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[801] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[802] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[803] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[804] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[805] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[806] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[807] = sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[808] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[809] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[810] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[811] = sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[812] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[813] = sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[814] = ~sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[815] = sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[816] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[817] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[818] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[819] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[820] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[821] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[822] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[823] = sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[824] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[825] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[826] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[827] = sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[828] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[829] = sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[830] = ~sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[831] = sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[832] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[833] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[834] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[835] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[836] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[837] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[838] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[839] = sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[840] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[841] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[842] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[843] = sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[844] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[845] = sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[846] = ~sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[847] = sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[848] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[849] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[850] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[851] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[852] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[853] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[854] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[855] = sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[856] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[857] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[858] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[859] = sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[860] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[861] = sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[862] = ~sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[863] = sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[864] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[865] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[866] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[867] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[868] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[869] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[870] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[871] = sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[872] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[873] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[874] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[875] = sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[876] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[877] = sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[878] = ~sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[879] = sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[880] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[881] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[882] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[883] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[884] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[885] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[886] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[887] = sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[888] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[889] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[890] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[891] = sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[892] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[893] = sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[894] = ~sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[895] = sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
	 address[896] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
	 address[897] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
	 address[898] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
	 address[899] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
	 address[900] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
	 address[901] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
	 address[902] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
	 address[903] = sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
	 address[904] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
	 address[905] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
	 address[906] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
	 address[907] = sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
	 address[908] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
	 address[909] = sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
	 address[910] = ~sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
	 address[911] = sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
	 address[912] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
	 address[913] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
	 address[914] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
	 address[915] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
	 address[916] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
	 address[917] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
	 address[918] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
	 address[919] = sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
	 address[920] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
	 address[921] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
	 address[922] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
	 address[923] = sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
	 address[924] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
	 address[925] = sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
	 address[926] = ~sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
	 address[927] = sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
	 address[928] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
	 address[929] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
	 address[930] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
	 address[931] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
	 address[932] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
	 address[933] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
	 address[934] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
	 address[935] = sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
	 address[936] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
	 address[937] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
	 address[938] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
	 address[939] = sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
	 address[940] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
	 address[941] = sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
	 address[942] = ~sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
	 address[943] = sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
	 address[944] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
	 address[945] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
	 address[946] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
	 address[947] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
	 address[948] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
	 address[949] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
	 address[950] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
	 address[951] = sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
	 address[952] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
	 address[953] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
	 address[954] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
	 address[955] = sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
	 address[956] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
	 address[957] = sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
	 address[958] = ~sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
	 address[959] = sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
	 address[960] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
	 address[961] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
	 address[962] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
	 address[963] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
	 address[964] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
	 address[965] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
	 address[966] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
	 address[967] = sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
	 address[968] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
	 address[969] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
	 address[970] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
	 address[971] = sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
	 address[972] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
	 address[973] = sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
	 address[974] = ~sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
	 address[975] = sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
	 address[976] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
	 address[977] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
	 address[978] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
	 address[979] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
	 address[980] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
	 address[981] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
	 address[982] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
	 address[983] = sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
	 address[984] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
	 address[985] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
	 address[986] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
	 address[987] = sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
	 address[988] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
	 address[989] = sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
	 address[990] = ~sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
	 address[991] = sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
	 address[992] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
	 address[993] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
	 address[994] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
	 address[995] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
	 address[996] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
	 address[997] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
	 address[998] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
	 address[999] = sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
	 address[1000] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
	 address[1001] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
	 address[1002] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
	 address[1003] = sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
	 address[1004] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
	 address[1005] = sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
	 address[1006] = ~sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
	 address[1007] = sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
	 address[1008] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
	 address[1009] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
	 address[1010] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
	 address[1011] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
	 address[1012] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
	 address[1013] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
	 address[1014] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
	 address[1015] = sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
	 address[1016] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
	 address[1017] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
	 address[1018] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
	 address[1019] = sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
	 address[1020] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
	 address[1021] = sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
	 address[1022] = ~sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
	 address[1023] = sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & sel[9];

    end

endmodule


`default_nettype wire
