module IMPACTSram (

`ifdef USE_POWER_PINS
    inout vccd1,	// User area 2 1.8v supply
    inout vssd1,	// User area 2 digital ground
`endif



//   inout vccd1, // User area 1 1.8V supply
//   inout vssd1, // User area 1 digital ground


    // Wishbone Slave ports (WB MI A)

    // Logic Analyzer Signals

    // IRQ
    input PRE,
    input ReadEn,
    input WriteEn,
    input [1023:0] Address,
    input [31:0] DataIn,
    output [31:0] DataOut

);

wire [1023:0] WL;
assign WL = Address;

//wire [31:0] WL_Bank01;
//################################################
//Creates the Four Word Decoders Instences for the Four Memory Banks
//################################################

//Bank01 SRAM Block
full_sram full_sram(
`ifdef USE_POWER_PINS
	.vccd1(vccd1),	// User area 1 1.8V power
	.vssd1(vssd1),	// User area 1 digital ground
`endif

.PRE(PRE),
.readen(ReadEn),
.writeen(WriteEn),

.DataIn0(DataIn [0]),
.DataIn1(DataIn [1]),
.DataIn2(DataIn [2]),
.DataIn3(DataIn [3]),
.DataIn4(DataIn [4]),
.DataIn5(DataIn [5]),
.DataIn6(DataIn [6]),
.DataIn7(DataIn [7]),
.DataIn8(DataIn [8]),
.DataIn9(DataIn [9]),
.DataIn10(DataIn [10]),
.DataIn11(DataIn [11]),
.DataIn12(DataIn [12]),
.DataIn13(DataIn [13]),
.DataIn14(DataIn [14]),
.DataIn15(DataIn [15]),
.DataIn16(DataIn [16]),
.DataIn17(DataIn [17]),
.DataIn18(DataIn [18]),
.DataIn19(DataIn [19]),
.DataIn20(DataIn [20]),
.DataIn21(DataIn [21]),
.DataIn22(DataIn [22]),
.DataIn23(DataIn [23]),
.DataIn24(DataIn [24]),
.DataIn25(DataIn [25]),
.DataIn26(DataIn [26]),
.DataIn27(DataIn [27]),
.DataIn28(DataIn [28]),
.DataIn29(DataIn [29]),
.DataIn30(DataIn [30]),
.DataIn31(DataIn [31]),


.DataOut0(DataOut [0]),
.DataOut1(DataOut [1]),
.DataOut2(DataOut [2]),
.DataOut3(DataOut [3]),
.DataOut4(DataOut [4]),
.DataOut5(DataOut [5]),
.DataOut6(DataOut [6]),
.DataOut7(DataOut [7]),
.DataOut8(DataOut [8]),
.DataOut9(DataOut [9]),
.DataOut10(DataOut [10]),
.DataOut11(DataOut [11]),
.DataOut12(DataOut [12]),
.DataOut13(DataOut [13]),
.DataOut14(DataOut [14]),
.DataOut15(DataOut [15]),
.DataOut16(DataOut [16]),
.DataOut17(DataOut [17]),
.DataOut18(DataOut [18]),
.DataOut19(DataOut [19]),
.DataOut20(DataOut [20]),
.DataOut21(DataOut [21]),
.DataOut22(DataOut [22]),
.DataOut23(DataOut [23]),
.DataOut24(DataOut [24]),
.DataOut25(DataOut [25]),
.DataOut26(DataOut [26]),
.DataOut27(DataOut [27]),
.DataOut28(DataOut [28]),
.DataOut29(DataOut [29]),
.DataOut30(DataOut [30]),
.DataOut31(DataOut [31]),


.WL0(WL [0]),
.WL1(WL [1]),
.WL2(WL [2]),
.WL3(WL [3]),
.WL4(WL [4]),
.WL5(WL [5]),
.WL6(WL [6]),
.WL7(WL [7]),
.WL8(WL [8]),
.WL9(WL [9]),
.WL10(WL [10]),
.WL11(WL [11]),
.WL12(WL [12]),
.WL13(WL [13]),
.WL14(WL [14]),
.WL15(WL [15]),
.WL16(WL [16]),
.WL17(WL [17]),
.WL18(WL [18]),
.WL19(WL [19]),
.WL20(WL [20]),
.WL21(WL [21]),
.WL22(WL [22]),
.WL23(WL [23]),
.WL24(WL [24]),
.WL25(WL [25]),
.WL26(WL [26]),
.WL27(WL [27]),
.WL28(WL [28]),
.WL29(WL [29]),
.WL30(WL [30]),
.WL31(WL [31]),
.WL32(WL [32]),
.WL33(WL [33]),
.WL34(WL [34]),
.WL35(WL [35]),
.WL36(WL [36]),
.WL37(WL [37]),
.WL38(WL [38]),
.WL39(WL [39]),
.WL40(WL [40]),
.WL41(WL [41]),
.WL42(WL [42]),
.WL43(WL [43]),
.WL44(WL [44]),
.WL45(WL [45]),
.WL46(WL [46]),
.WL47(WL [47]),
.WL48(WL [48]),
.WL49(WL [49]),
.WL50(WL [50]),
.WL51(WL [51]),
.WL52(WL [52]),
.WL53(WL [53]),
.WL54(WL [54]),
.WL55(WL [55]),
.WL56(WL [56]),
.WL57(WL [57]),
.WL58(WL [58]),
.WL59(WL [59]),
.WL60(WL [60]),
.WL61(WL [61]),
.WL62(WL [62]),
.WL63(WL [63]),
.WL64(WL [64]),
.WL65(WL [65]),
.WL66(WL [66]),
.WL67(WL [67]),
.WL68(WL [68]),
.WL69(WL [69]),
.WL70(WL [70]),
.WL71(WL [71]),
.WL72(WL [72]),
.WL73(WL [73]),
.WL74(WL [74]),
.WL75(WL [75]),
.WL76(WL [76]),
.WL77(WL [77]),
.WL78(WL [78]),
.WL79(WL [79]),
.WL80(WL [80]),
.WL81(WL [81]),
.WL82(WL [82]),
.WL83(WL [83]),
.WL84(WL [84]),
.WL85(WL [85]),
.WL86(WL [86]),
.WL87(WL [87]),
.WL88(WL [88]),
.WL89(WL [89]),
.WL90(WL [90]),
.WL91(WL [91]),
.WL92(WL [92]),
.WL93(WL [93]),
.WL94(WL [94]),
.WL95(WL [95]),
.WL96(WL [96]),
.WL97(WL [97]),
.WL98(WL [98]),
.WL99(WL [99]),
.WL100(WL [100]),
.WL101(WL [101]),
.WL102(WL [102]),
.WL103(WL [103]),
.WL104(WL [104]),
.WL105(WL [105]),
.WL106(WL [106]),
.WL107(WL [107]),
.WL108(WL [108]),
.WL109(WL [109]),
.WL110(WL [110]),
.WL111(WL [111]),
.WL112(WL [112]),
.WL113(WL [113]),
.WL114(WL [114]),
.WL115(WL [115]),
.WL116(WL [116]),
.WL117(WL [117]),
.WL118(WL [118]),
.WL119(WL [119]),
.WL120(WL [120]),
.WL121(WL [121]),
.WL122(WL [122]),
.WL123(WL [123]),
.WL124(WL [124]),
.WL125(WL [125]),
.WL126(WL [126]),
.WL127(WL [127]),
.WL128(WL [128]),
.WL129(WL [129]),
.WL130(WL [130]),
.WL131(WL [131]),
.WL132(WL [132]),
.WL133(WL [133]),
.WL134(WL [134]),
.WL135(WL [135]),
.WL136(WL [136]),
.WL137(WL [137]),
.WL138(WL [138]),
.WL139(WL [139]),
.WL140(WL [140]),
.WL141(WL [141]),
.WL142(WL [142]),
.WL143(WL [143]),
.WL144(WL [144]),
.WL145(WL [145]),
.WL146(WL [146]),
.WL147(WL [147]),
.WL148(WL [148]),
.WL149(WL [149]),
.WL150(WL [150]),
.WL151(WL [151]),
.WL152(WL [152]),
.WL153(WL [153]),
.WL154(WL [154]),
.WL155(WL [155]),
.WL156(WL [156]),
.WL157(WL [157]),
.WL158(WL [158]),
.WL159(WL [159]),
.WL160(WL [160]),
.WL161(WL [161]),
.WL162(WL [162]),
.WL163(WL [163]),
.WL164(WL [164]),
.WL165(WL [165]),
.WL166(WL [166]),
.WL167(WL [167]),
.WL168(WL [168]),
.WL169(WL [169]),
.WL170(WL [170]),
.WL171(WL [171]),
.WL172(WL [172]),
.WL173(WL [173]),
.WL174(WL [174]),
.WL175(WL [175]),
.WL176(WL [176]),
.WL177(WL [177]),
.WL178(WL [178]),
.WL179(WL [179]),
.WL180(WL [180]),
.WL181(WL [181]),
.WL182(WL [182]),
.WL183(WL [183]),
.WL184(WL [184]),
.WL185(WL [185]),
.WL186(WL [186]),
.WL187(WL [187]),
.WL188(WL [188]),
.WL189(WL [189]),
.WL190(WL [190]),
.WL191(WL [191]),
.WL192(WL [192]),
.WL193(WL [193]),
.WL194(WL [194]),
.WL195(WL [195]),
.WL196(WL [196]),
.WL197(WL [197]),
.WL198(WL [198]),
.WL199(WL [199]),
.WL200(WL [200]),
.WL201(WL [201]),
.WL202(WL [202]),
.WL203(WL [203]),
.WL204(WL [204]),
.WL205(WL [205]),
.WL206(WL [206]),
.WL207(WL [207]),
.WL208(WL [208]),
.WL209(WL [209]),
.WL210(WL [210]),
.WL211(WL [211]),
.WL212(WL [212]),
.WL213(WL [213]),
.WL214(WL [214]),
.WL215(WL [215]),
.WL216(WL [216]),
.WL217(WL [217]),
.WL218(WL [218]),
.WL219(WL [219]),
.WL220(WL [220]),
.WL221(WL [221]),
.WL222(WL [222]),
.WL223(WL [223]),
.WL224(WL [224]),
.WL225(WL [225]),
.WL226(WL [226]),
.WL227(WL [227]),
.WL228(WL [228]),
.WL229(WL [229]),
.WL230(WL [230]),
.WL231(WL [231]),
.WL232(WL [232]),
.WL233(WL [233]),
.WL234(WL [234]),
.WL235(WL [235]),
.WL236(WL [236]),
.WL237(WL [237]),
.WL238(WL [238]),
.WL239(WL [239]),
.WL240(WL [240]),
.WL241(WL [241]),
.WL242(WL [242]),
.WL243(WL [243]),
.WL244(WL [244]),
.WL245(WL [245]),
.WL246(WL [246]),
.WL247(WL [247]),
.WL248(WL [248]),
.WL249(WL [249]),
.WL250(WL [250]),
.WL251(WL [251]),
.WL252(WL [252]),
.WL253(WL [253]),
.WL254(WL [254]),
.WL255(WL [255]),
.WL256(WL [256]),
.WL257(WL [257]),
.WL258(WL [258]),
.WL259(WL [259]),
.WL260(WL [260]),
.WL261(WL [261]),
.WL262(WL [262]),
.WL263(WL [263]),
.WL264(WL [264]),
.WL265(WL [265]),
.WL266(WL [266]),
.WL267(WL [267]),
.WL268(WL [268]),
.WL269(WL [269]),
.WL270(WL [270]),
.WL271(WL [271]),
.WL272(WL [272]),
.WL273(WL [273]),
.WL274(WL [274]),
.WL275(WL [275]),
.WL276(WL [276]),
.WL277(WL [277]),
.WL278(WL [278]),
.WL279(WL [279]),
.WL280(WL [280]),
.WL281(WL [281]),
.WL282(WL [282]),
.WL283(WL [283]),
.WL284(WL [284]),
.WL285(WL [285]),
.WL286(WL [286]),
.WL287(WL [287]),
.WL288(WL [288]),
.WL289(WL [289]),
.WL290(WL [290]),
.WL291(WL [291]),
.WL292(WL [292]),
.WL293(WL [293]),
.WL294(WL [294]),
.WL295(WL [295]),
.WL296(WL [296]),
.WL297(WL [297]),
.WL298(WL [298]),
.WL299(WL [299]),
.WL300(WL [300]),
.WL301(WL [301]),
.WL302(WL [302]),
.WL303(WL [303]),
.WL304(WL [304]),
.WL305(WL [305]),
.WL306(WL [306]),
.WL307(WL [307]),
.WL308(WL [308]),
.WL309(WL [309]),
.WL310(WL [310]),
.WL311(WL [311]),
.WL312(WL [312]),
.WL313(WL [313]),
.WL314(WL [314]),
.WL315(WL [315]),
.WL316(WL [316]),
.WL317(WL [317]),
.WL318(WL [318]),
.WL319(WL [319]),
.WL320(WL [320]),
.WL321(WL [321]),
.WL322(WL [322]),
.WL323(WL [323]),
.WL324(WL [324]),
.WL325(WL [325]),
.WL326(WL [326]),
.WL327(WL [327]),
.WL328(WL [328]),
.WL329(WL [329]),
.WL330(WL [330]),
.WL331(WL [331]),
.WL332(WL [332]),
.WL333(WL [333]),
.WL334(WL [334]),
.WL335(WL [335]),
.WL336(WL [336]),
.WL337(WL [337]),
.WL338(WL [338]),
.WL339(WL [339]),
.WL340(WL [340]),
.WL341(WL [341]),
.WL342(WL [342]),
.WL343(WL [343]),
.WL344(WL [344]),
.WL345(WL [345]),
.WL346(WL [346]),
.WL347(WL [347]),
.WL348(WL [348]),
.WL349(WL [349]),
.WL350(WL [350]),
.WL351(WL [351]),
.WL352(WL [352]),
.WL353(WL [353]),
.WL354(WL [354]),
.WL355(WL [355]),
.WL356(WL [356]),
.WL357(WL [357]),
.WL358(WL [358]),
.WL359(WL [359]),
.WL360(WL [360]),
.WL361(WL [361]),
.WL362(WL [362]),
.WL363(WL [363]),
.WL364(WL [364]),
.WL365(WL [365]),
.WL366(WL [366]),
.WL367(WL [367]),
.WL368(WL [368]),
.WL369(WL [369]),
.WL370(WL [370]),
.WL371(WL [371]),
.WL372(WL [372]),
.WL373(WL [373]),
.WL374(WL [374]),
.WL375(WL [375]),
.WL376(WL [376]),
.WL377(WL [377]),
.WL378(WL [378]),
.WL379(WL [379]),
.WL380(WL [380]),
.WL381(WL [381]),
.WL382(WL [382]),
.WL383(WL [383]),
.WL384(WL [384]),
.WL385(WL [385]),
.WL386(WL [386]),
.WL387(WL [387]),
.WL388(WL [388]),
.WL389(WL [389]),
.WL390(WL [390]),
.WL391(WL [391]),
.WL392(WL [392]),
.WL393(WL [393]),
.WL394(WL [394]),
.WL395(WL [395]),
.WL396(WL [396]),
.WL397(WL [397]),
.WL398(WL [398]),
.WL399(WL [399]),
.WL400(WL [400]),
.WL401(WL [401]),
.WL402(WL [402]),
.WL403(WL [403]),
.WL404(WL [404]),
.WL405(WL [405]),
.WL406(WL [406]),
.WL407(WL [407]),
.WL408(WL [408]),
.WL409(WL [409]),
.WL410(WL [410]),
.WL411(WL [411]),
.WL412(WL [412]),
.WL413(WL [413]),
.WL414(WL [414]),
.WL415(WL [415]),
.WL416(WL [416]),
.WL417(WL [417]),
.WL418(WL [418]),
.WL419(WL [419]),
.WL420(WL [420]),
.WL421(WL [421]),
.WL422(WL [422]),
.WL423(WL [423]),
.WL424(WL [424]),
.WL425(WL [425]),
.WL426(WL [426]),
.WL427(WL [427]),
.WL428(WL [428]),
.WL429(WL [429]),
.WL430(WL [430]),
.WL431(WL [431]),
.WL432(WL [432]),
.WL433(WL [433]),
.WL434(WL [434]),
.WL435(WL [435]),
.WL436(WL [436]),
.WL437(WL [437]),
.WL438(WL [438]),
.WL439(WL [439]),
.WL440(WL [440]),
.WL441(WL [441]),
.WL442(WL [442]),
.WL443(WL [443]),
.WL444(WL [444]),
.WL445(WL [445]),
.WL446(WL [446]),
.WL447(WL [447]),
.WL448(WL [448]),
.WL449(WL [449]),
.WL450(WL [450]),
.WL451(WL [451]),
.WL452(WL [452]),
.WL453(WL [453]),
.WL454(WL [454]),
.WL455(WL [455]),
.WL456(WL [456]),
.WL457(WL [457]),
.WL458(WL [458]),
.WL459(WL [459]),
.WL460(WL [460]),
.WL461(WL [461]),
.WL462(WL [462]),
.WL463(WL [463]),
.WL464(WL [464]),
.WL465(WL [465]),
.WL466(WL [466]),
.WL467(WL [467]),
.WL468(WL [468]),
.WL469(WL [469]),
.WL470(WL [470]),
.WL471(WL [471]),
.WL472(WL [472]),
.WL473(WL [473]),
.WL474(WL [474]),
.WL475(WL [475]),
.WL476(WL [476]),
.WL477(WL [477]),
.WL478(WL [478]),
.WL479(WL [479]),
.WL480(WL [480]),
.WL481(WL [481]),
.WL482(WL [482]),
.WL483(WL [483]),
.WL484(WL [484]),
.WL485(WL [485]),
.WL486(WL [486]),
.WL487(WL [487]),
.WL488(WL [488]),
.WL489(WL [489]),
.WL490(WL [490]),
.WL491(WL [491]),
.WL492(WL [492]),
.WL493(WL [493]),
.WL494(WL [494]),
.WL495(WL [495]),
.WL496(WL [496]),
.WL497(WL [497]),
.WL498(WL [498]),
.WL499(WL [499]),
.WL500(WL [500]),
.WL501(WL [501]),
.WL502(WL [502]),
.WL503(WL [503]),
.WL504(WL [504]),
.WL505(WL [505]),
.WL506(WL [506]),
.WL507(WL [507]),
.WL508(WL [508]),
.WL509(WL [509]),
.WL510(WL [510]),
.WL511(WL [511]),
.WL512(WL [512]),
.WL513(WL [513]),
.WL514(WL [514]),
.WL515(WL [515]),
.WL516(WL [516]),
.WL517(WL [517]),
.WL518(WL [518]),
.WL519(WL [519]),
.WL520(WL [520]),
.WL521(WL [521]),
.WL522(WL [522]),
.WL523(WL [523]),
.WL524(WL [524]),
.WL525(WL [525]),
.WL526(WL [526]),
.WL527(WL [527]),
.WL528(WL [528]),
.WL529(WL [529]),
.WL530(WL [530]),
.WL531(WL [531]),
.WL532(WL [532]),
.WL533(WL [533]),
.WL534(WL [534]),
.WL535(WL [535]),
.WL536(WL [536]),
.WL537(WL [537]),
.WL538(WL [538]),
.WL539(WL [539]),
.WL540(WL [540]),
.WL541(WL [541]),
.WL542(WL [542]),
.WL543(WL [543]),
.WL544(WL [544]),
.WL545(WL [545]),
.WL546(WL [546]),
.WL547(WL [547]),
.WL548(WL [548]),
.WL549(WL [549]),
.WL550(WL [550]),
.WL551(WL [551]),
.WL552(WL [552]),
.WL553(WL [553]),
.WL554(WL [554]),
.WL555(WL [555]),
.WL556(WL [556]),
.WL557(WL [557]),
.WL558(WL [558]),
.WL559(WL [559]),
.WL560(WL [560]),
.WL561(WL [561]),
.WL562(WL [562]),
.WL563(WL [563]),
.WL564(WL [564]),
.WL565(WL [565]),
.WL566(WL [566]),
.WL567(WL [567]),
.WL568(WL [568]),
.WL569(WL [569]),
.WL570(WL [570]),
.WL571(WL [571]),
.WL572(WL [572]),
.WL573(WL [573]),
.WL574(WL [574]),
.WL575(WL [575]),
.WL576(WL [576]),
.WL577(WL [577]),
.WL578(WL [578]),
.WL579(WL [579]),
.WL580(WL [580]),
.WL581(WL [581]),
.WL582(WL [582]),
.WL583(WL [583]),
.WL584(WL [584]),
.WL585(WL [585]),
.WL586(WL [586]),
.WL587(WL [587]),
.WL588(WL [588]),
.WL589(WL [589]),
.WL590(WL [590]),
.WL591(WL [591]),
.WL592(WL [592]),
.WL593(WL [593]),
.WL594(WL [594]),
.WL595(WL [595]),
.WL596(WL [596]),
.WL597(WL [597]),
.WL598(WL [598]),
.WL599(WL [599]),
.WL600(WL [600]),
.WL601(WL [601]),
.WL602(WL [602]),
.WL603(WL [603]),
.WL604(WL [604]),
.WL605(WL [605]),
.WL606(WL [606]),
.WL607(WL [607]),
.WL608(WL [608]),
.WL609(WL [609]),
.WL610(WL [610]),
.WL611(WL [611]),
.WL612(WL [612]),
.WL613(WL [613]),
.WL614(WL [614]),
.WL615(WL [615]),
.WL616(WL [616]),
.WL617(WL [617]),
.WL618(WL [618]),
.WL619(WL [619]),
.WL620(WL [620]),
.WL621(WL [621]),
.WL622(WL [622]),
.WL623(WL [623]),
.WL624(WL [624]),
.WL625(WL [625]),
.WL626(WL [626]),
.WL627(WL [627]),
.WL628(WL [628]),
.WL629(WL [629]),
.WL630(WL [630]),
.WL631(WL [631]),
.WL632(WL [632]),
.WL633(WL [633]),
.WL634(WL [634]),
.WL635(WL [635]),
.WL636(WL [636]),
.WL637(WL [637]),
.WL638(WL [638]),
.WL639(WL [639]),
.WL640(WL [640]),
.WL641(WL [641]),
.WL642(WL [642]),
.WL643(WL [643]),
.WL644(WL [644]),
.WL645(WL [645]),
.WL646(WL [646]),
.WL647(WL [647]),
.WL648(WL [648]),
.WL649(WL [649]),
.WL650(WL [650]),
.WL651(WL [651]),
.WL652(WL [652]),
.WL653(WL [653]),
.WL654(WL [654]),
.WL655(WL [655]),
.WL656(WL [656]),
.WL657(WL [657]),
.WL658(WL [658]),
.WL659(WL [659]),
.WL660(WL [660]),
.WL661(WL [661]),
.WL662(WL [662]),
.WL663(WL [663]),
.WL664(WL [664]),
.WL665(WL [665]),
.WL666(WL [666]),
.WL667(WL [667]),
.WL668(WL [668]),
.WL669(WL [669]),
.WL670(WL [670]),
.WL671(WL [671]),
.WL672(WL [672]),
.WL673(WL [673]),
.WL674(WL [674]),
.WL675(WL [675]),
.WL676(WL [676]),
.WL677(WL [677]),
.WL678(WL [678]),
.WL679(WL [679]),
.WL680(WL [680]),
.WL681(WL [681]),
.WL682(WL [682]),
.WL683(WL [683]),
.WL684(WL [684]),
.WL685(WL [685]),
.WL686(WL [686]),
.WL687(WL [687]),
.WL688(WL [688]),
.WL689(WL [689]),
.WL690(WL [690]),
.WL691(WL [691]),
.WL692(WL [692]),
.WL693(WL [693]),
.WL694(WL [694]),
.WL695(WL [695]),
.WL696(WL [696]),
.WL697(WL [697]),
.WL698(WL [698]),
.WL699(WL [699]),
.WL700(WL [700]),
.WL701(WL [701]),
.WL702(WL [702]),
.WL703(WL [703]),
.WL704(WL [704]),
.WL705(WL [705]),
.WL706(WL [706]),
.WL707(WL [707]),
.WL708(WL [708]),
.WL709(WL [709]),
.WL710(WL [710]),
.WL711(WL [711]),
.WL712(WL [712]),
.WL713(WL [713]),
.WL714(WL [714]),
.WL715(WL [715]),
.WL716(WL [716]),
.WL717(WL [717]),
.WL718(WL [718]),
.WL719(WL [719]),
.WL720(WL [720]),
.WL721(WL [721]),
.WL722(WL [722]),
.WL723(WL [723]),
.WL724(WL [724]),
.WL725(WL [725]),
.WL726(WL [726]),
.WL727(WL [727]),
.WL728(WL [728]),
.WL729(WL [729]),
.WL730(WL [730]),
.WL731(WL [731]),
.WL732(WL [732]),
.WL733(WL [733]),
.WL734(WL [734]),
.WL735(WL [735]),
.WL736(WL [736]),
.WL737(WL [737]),
.WL738(WL [738]),
.WL739(WL [739]),
.WL740(WL [740]),
.WL741(WL [741]),
.WL742(WL [742]),
.WL743(WL [743]),
.WL744(WL [744]),
.WL745(WL [745]),
.WL746(WL [746]),
.WL747(WL [747]),
.WL748(WL [748]),
.WL749(WL [749]),
.WL750(WL [750]),
.WL751(WL [751]),
.WL752(WL [752]),
.WL753(WL [753]),
.WL754(WL [754]),
.WL755(WL [755]),
.WL756(WL [756]),
.WL757(WL [757]),
.WL758(WL [758]),
.WL759(WL [759]),
.WL760(WL [760]),
.WL761(WL [761]),
.WL762(WL [762]),
.WL763(WL [763]),
.WL764(WL [764]),
.WL765(WL [765]),
.WL766(WL [766]),
.WL767(WL [767]),
.WL768(WL [768]),
.WL769(WL [769]),
.WL770(WL [770]),
.WL771(WL [771]),
.WL772(WL [772]),
.WL773(WL [773]),
.WL774(WL [774]),
.WL775(WL [775]),
.WL776(WL [776]),
.WL777(WL [777]),
.WL778(WL [778]),
.WL779(WL [779]),
.WL780(WL [780]),
.WL781(WL [781]),
.WL782(WL [782]),
.WL783(WL [783]),
.WL784(WL [784]),
.WL785(WL [785]),
.WL786(WL [786]),
.WL787(WL [787]),
.WL788(WL [788]),
.WL789(WL [789]),
.WL790(WL [790]),
.WL791(WL [791]),
.WL792(WL [792]),
.WL793(WL [793]),
.WL794(WL [794]),
.WL795(WL [795]),
.WL796(WL [796]),
.WL797(WL [797]),
.WL798(WL [798]),
.WL799(WL [799]),
.WL800(WL [800]),
.WL801(WL [801]),
.WL802(WL [802]),
.WL803(WL [803]),
.WL804(WL [804]),
.WL805(WL [805]),
.WL806(WL [806]),
.WL807(WL [807]),
.WL808(WL [808]),
.WL809(WL [809]),
.WL810(WL [810]),
.WL811(WL [811]),
.WL812(WL [812]),
.WL813(WL [813]),
.WL814(WL [814]),
.WL815(WL [815]),
.WL816(WL [816]),
.WL817(WL [817]),
.WL818(WL [818]),
.WL819(WL [819]),
.WL820(WL [820]),
.WL821(WL [821]),
.WL822(WL [822]),
.WL823(WL [823]),
.WL824(WL [824]),
.WL825(WL [825]),
.WL826(WL [826]),
.WL827(WL [827]),
.WL828(WL [828]),
.WL829(WL [829]),
.WL830(WL [830]),
.WL831(WL [831]),
.WL832(WL [832]),
.WL833(WL [833]),
.WL834(WL [834]),
.WL835(WL [835]),
.WL836(WL [836]),
.WL837(WL [837]),
.WL838(WL [838]),
.WL839(WL [839]),
.WL840(WL [840]),
.WL841(WL [841]),
.WL842(WL [842]),
.WL843(WL [843]),
.WL844(WL [844]),
.WL845(WL [845]),
.WL846(WL [846]),
.WL847(WL [847]),
.WL848(WL [848]),
.WL849(WL [849]),
.WL850(WL [850]),
.WL851(WL [851]),
.WL852(WL [852]),
.WL853(WL [853]),
.WL854(WL [854]),
.WL855(WL [855]),
.WL856(WL [856]),
.WL857(WL [857]),
.WL858(WL [858]),
.WL859(WL [859]),
.WL860(WL [860]),
.WL861(WL [861]),
.WL862(WL [862]),
.WL863(WL [863]),
.WL864(WL [864]),
.WL865(WL [865]),
.WL866(WL [866]),
.WL867(WL [867]),
.WL868(WL [868]),
.WL869(WL [869]),
.WL870(WL [870]),
.WL871(WL [871]),
.WL872(WL [872]),
.WL873(WL [873]),
.WL874(WL [874]),
.WL875(WL [875]),
.WL876(WL [876]),
.WL877(WL [877]),
.WL878(WL [878]),
.WL879(WL [879]),
.WL880(WL [880]),
.WL881(WL [881]),
.WL882(WL [882]),
.WL883(WL [883]),
.WL884(WL [884]),
.WL885(WL [885]),
.WL886(WL [886]),
.WL887(WL [887]),
.WL888(WL [888]),
.WL889(WL [889]),
.WL890(WL [890]),
.WL891(WL [891]),
.WL892(WL [892]),
.WL893(WL [893]),
.WL894(WL [894]),
.WL895(WL [895]),
.WL896(WL [896]),
.WL897(WL [897]),
.WL898(WL [898]),
.WL899(WL [899]),
.WL900(WL [900]),
.WL901(WL [901]),
.WL902(WL [902]),
.WL903(WL [903]),
.WL904(WL [904]),
.WL905(WL [905]),
.WL906(WL [906]),
.WL907(WL [907]),
.WL908(WL [908]),
.WL909(WL [909]),
.WL910(WL [910]),
.WL911(WL [911]),
.WL912(WL [912]),
.WL913(WL [913]),
.WL914(WL [914]),
.WL915(WL [915]),
.WL916(WL [916]),
.WL917(WL [917]),
.WL918(WL [918]),
.WL919(WL [919]),
.WL920(WL [920]),
.WL921(WL [921]),
.WL922(WL [922]),
.WL923(WL [923]),
.WL924(WL [924]),
.WL925(WL [925]),
.WL926(WL [926]),
.WL927(WL [927]),
.WL928(WL [928]),
.WL929(WL [929]),
.WL930(WL [930]),
.WL931(WL [931]),
.WL932(WL [932]),
.WL933(WL [933]),
.WL934(WL [934]),
.WL935(WL [935]),
.WL936(WL [936]),
.WL937(WL [937]),
.WL938(WL [938]),
.WL939(WL [939]),
.WL940(WL [940]),
.WL941(WL [941]),
.WL942(WL [942]),
.WL943(WL [943]),
.WL944(WL [944]),
.WL945(WL [945]),
.WL946(WL [946]),
.WL947(WL [947]),
.WL948(WL [948]),
.WL949(WL [949]),
.WL950(WL [950]),
.WL951(WL [951]),
.WL952(WL [952]),
.WL953(WL [953]),
.WL954(WL [954]),
.WL955(WL [955]),
.WL956(WL [956]),
.WL957(WL [957]),
.WL958(WL [958]),
.WL959(WL [959]),
.WL960(WL [960]),
.WL961(WL [961]),
.WL962(WL [962]),
.WL963(WL [963]),
.WL964(WL [964]),
.WL965(WL [965]),
.WL966(WL [966]),
.WL967(WL [967]),
.WL968(WL [968]),
.WL969(WL [969]),
.WL970(WL [970]),
.WL971(WL [971]),
.WL972(WL [972]),
.WL973(WL [973]),
.WL974(WL [974]),
.WL975(WL [975]),
.WL976(WL [976]),
.WL977(WL [977]),
.WL978(WL [978]),
.WL979(WL [979]),
.WL980(WL [980]),
.WL981(WL [981]),
.WL982(WL [982]),
.WL983(WL [983]),
.WL984(WL [984]),
.WL985(WL [985]),
.WL986(WL [986]),
.WL987(WL [987]),
.WL988(WL [988]),
.WL989(WL [989]),
.WL990(WL [990]),
.WL991(WL [991]),
.WL992(WL [992]),
.WL993(WL [993]),
.WL994(WL [994]),
.WL995(WL [995]),
.WL996(WL [996]),
.WL997(WL [997]),
.WL998(WL [998]),
.WL999(WL [999]),
.WL1000(WL [1000]),
.WL1001(WL [1001]),
.WL1002(WL [1002]),
.WL1003(WL [1003]),
.WL1004(WL [1004]),
.WL1005(WL [1005]),
.WL1006(WL [1006]),
.WL1007(WL [1007]),
.WL1008(WL [1008]),
.WL1009(WL [1009]),
.WL1010(WL [1010]),
.WL1011(WL [1011]),
.WL1012(WL [1012]),
.WL1013(WL [1013]),
.WL1014(WL [1014]),
.WL1015(WL [1015]),
.WL1016(WL [1016]),
.WL1017(WL [1017]),
.WL1018(WL [1018]),
.WL1019(WL [1019]),
.WL1020(WL [1020]),
.WL1021(WL [1021]),
.WL1022(WL [1022]),
.WL1023(WL [1023])

);

endmodule

(* blackbox *)
module full_sram (

`ifdef USE_POWER_PINS
	inout vccd1,	// User area 1 1.8V power
	inout vssd1,	// User area 1 digital ground
`endif

input PRE,
input readen,
input writeen,

input DataIn0,
input DataIn1,
input DataIn2,
input DataIn3,
input DataIn4,
input DataIn5,
input DataIn6,
input DataIn7,
input DataIn8,
input DataIn9,
input DataIn10,
input DataIn11,
input DataIn12,
input DataIn13,
input DataIn14,
input DataIn15,
input DataIn16,
input DataIn17,
input DataIn18,
input DataIn19,
input DataIn20,
input DataIn21,
input DataIn22,
input DataIn23,
input DataIn24,
input DataIn25,
input DataIn26,
input DataIn27,
input DataIn28,
input DataIn29,
input DataIn30,
input DataIn31,

output DataOut0,
output DataOut1,
output DataOut2,
output DataOut3,
output DataOut4,
output DataOut5,
output DataOut6,
output DataOut7,
output DataOut8,
output DataOut9,
output DataOut10,
output DataOut11,
output DataOut12,
output DataOut13,
output DataOut14,
output DataOut15,
output DataOut16,
output DataOut17,
output DataOut18,
output DataOut19,
output DataOut20,
output DataOut21,
output DataOut22,
output DataOut23,
output DataOut24,
output DataOut25,
output DataOut26,
output DataOut27,
output DataOut28,
output DataOut29,
output DataOut30,
output DataOut31,

input WL0,
input WL1,
input WL2,
input WL3,
input WL4,
input WL5,
input WL6,
input WL7,
input WL8,
input WL9,
input WL10,
input WL11,
input WL12,
input WL13,
input WL14,
input WL15,
input WL16,
input WL17,
input WL18,
input WL19,
input WL20,
input WL21,
input WL22,
input WL23,
input WL24,
input WL25,
input WL26,
input WL27,
input WL28,
input WL29,
input WL30,
input WL31,
input WL32,
input WL33,
input WL34,
input WL35,
input WL36,
input WL37,
input WL38,
input WL39,
input WL40,
input WL41,
input WL42,
input WL43,
input WL44,
input WL45,
input WL46,
input WL47,
input WL48,
input WL49,
input WL50,
input WL51,
input WL52,
input WL53,
input WL54,
input WL55,
input WL56,
input WL57,
input WL58,
input WL59,
input WL60,
input WL61,
input WL62,
input WL63,
input WL64,
input WL65,
input WL66,
input WL67,
input WL68,
input WL69,
input WL70,
input WL71,
input WL72,
input WL73,
input WL74,
input WL75,
input WL76,
input WL77,
input WL78,
input WL79,
input WL80,
input WL81,
input WL82,
input WL83,
input WL84,
input WL85,
input WL86,
input WL87,
input WL88,
input WL89,
input WL90,
input WL91,
input WL92,
input WL93,
input WL94,
input WL95,
input WL96,
input WL97,
input WL98,
input WL99,
input WL100,
input WL101,
input WL102,
input WL103,
input WL104,
input WL105,
input WL106,
input WL107,
input WL108,
input WL109,
input WL110,
input WL111,
input WL112,
input WL113,
input WL114,
input WL115,
input WL116,
input WL117,
input WL118,
input WL119,
input WL120,
input WL121,
input WL122,
input WL123,
input WL124,
input WL125,
input WL126,
input WL127,
input WL128,
input WL129,
input WL130,
input WL131,
input WL132,
input WL133,
input WL134,
input WL135,
input WL136,
input WL137,
input WL138,
input WL139,
input WL140,
input WL141,
input WL142,
input WL143,
input WL144,
input WL145,
input WL146,
input WL147,
input WL148,
input WL149,
input WL150,
input WL151,
input WL152,
input WL153,
input WL154,
input WL155,
input WL156,
input WL157,
input WL158,
input WL159,
input WL160,
input WL161,
input WL162,
input WL163,
input WL164,
input WL165,
input WL166,
input WL167,
input WL168,
input WL169,
input WL170,
input WL171,
input WL172,
input WL173,
input WL174,
input WL175,
input WL176,
input WL177,
input WL178,
input WL179,
input WL180,
input WL181,
input WL182,
input WL183,
input WL184,
input WL185,
input WL186,
input WL187,
input WL188,
input WL189,
input WL190,
input WL191,
input WL192,
input WL193,
input WL194,
input WL195,
input WL196,
input WL197,
input WL198,
input WL199,
input WL200,
input WL201,
input WL202,
input WL203,
input WL204,
input WL205,
input WL206,
input WL207,
input WL208,
input WL209,
input WL210,
input WL211,
input WL212,
input WL213,
input WL214,
input WL215,
input WL216,
input WL217,
input WL218,
input WL219,
input WL220,
input WL221,
input WL222,
input WL223,
input WL224,
input WL225,
input WL226,
input WL227,
input WL228,
input WL229,
input WL230,
input WL231,
input WL232,
input WL233,
input WL234,
input WL235,
input WL236,
input WL237,
input WL238,
input WL239,
input WL240,
input WL241,
input WL242,
input WL243,
input WL244,
input WL245,
input WL246,
input WL247,
input WL248,
input WL249,
input WL250,
input WL251,
input WL252,
input WL253,
input WL254,
input WL255,
input WL256,
input WL257,
input WL258,
input WL259,
input WL260,
input WL261,
input WL262,
input WL263,
input WL264,
input WL265,
input WL266,
input WL267,
input WL268,
input WL269,
input WL270,
input WL271,
input WL272,
input WL273,
input WL274,
input WL275,
input WL276,
input WL277,
input WL278,
input WL279,
input WL280,
input WL281,
input WL282,
input WL283,
input WL284,
input WL285,
input WL286,
input WL287,
input WL288,
input WL289,
input WL290,
input WL291,
input WL292,
input WL293,
input WL294,
input WL295,
input WL296,
input WL297,
input WL298,
input WL299,
input WL300,
input WL301,
input WL302,
input WL303,
input WL304,
input WL305,
input WL306,
input WL307,
input WL308,
input WL309,
input WL310,
input WL311,
input WL312,
input WL313,
input WL314,
input WL315,
input WL316,
input WL317,
input WL318,
input WL319,
input WL320,
input WL321,
input WL322,
input WL323,
input WL324,
input WL325,
input WL326,
input WL327,
input WL328,
input WL329,
input WL330,
input WL331,
input WL332,
input WL333,
input WL334,
input WL335,
input WL336,
input WL337,
input WL338,
input WL339,
input WL340,
input WL341,
input WL342,
input WL343,
input WL344,
input WL345,
input WL346,
input WL347,
input WL348,
input WL349,
input WL350,
input WL351,
input WL352,
input WL353,
input WL354,
input WL355,
input WL356,
input WL357,
input WL358,
input WL359,
input WL360,
input WL361,
input WL362,
input WL363,
input WL364,
input WL365,
input WL366,
input WL367,
input WL368,
input WL369,
input WL370,
input WL371,
input WL372,
input WL373,
input WL374,
input WL375,
input WL376,
input WL377,
input WL378,
input WL379,
input WL380,
input WL381,
input WL382,
input WL383,
input WL384,
input WL385,
input WL386,
input WL387,
input WL388,
input WL389,
input WL390,
input WL391,
input WL392,
input WL393,
input WL394,
input WL395,
input WL396,
input WL397,
input WL398,
input WL399,
input WL400,
input WL401,
input WL402,
input WL403,
input WL404,
input WL405,
input WL406,
input WL407,
input WL408,
input WL409,
input WL410,
input WL411,
input WL412,
input WL413,
input WL414,
input WL415,
input WL416,
input WL417,
input WL418,
input WL419,
input WL420,
input WL421,
input WL422,
input WL423,
input WL424,
input WL425,
input WL426,
input WL427,
input WL428,
input WL429,
input WL430,
input WL431,
input WL432,
input WL433,
input WL434,
input WL435,
input WL436,
input WL437,
input WL438,
input WL439,
input WL440,
input WL441,
input WL442,
input WL443,
input WL444,
input WL445,
input WL446,
input WL447,
input WL448,
input WL449,
input WL450,
input WL451,
input WL452,
input WL453,
input WL454,
input WL455,
input WL456,
input WL457,
input WL458,
input WL459,
input WL460,
input WL461,
input WL462,
input WL463,
input WL464,
input WL465,
input WL466,
input WL467,
input WL468,
input WL469,
input WL470,
input WL471,
input WL472,
input WL473,
input WL474,
input WL475,
input WL476,
input WL477,
input WL478,
input WL479,
input WL480,
input WL481,
input WL482,
input WL483,
input WL484,
input WL485,
input WL486,
input WL487,
input WL488,
input WL489,
input WL490,
input WL491,
input WL492,
input WL493,
input WL494,
input WL495,
input WL496,
input WL497,
input WL498,
input WL499,
input WL500,
input WL501,
input WL502,
input WL503,
input WL504,
input WL505,
input WL506,
input WL507,
input WL508,
input WL509,
input WL510,
input WL511,
input WL512,
input WL513,
input WL514,
input WL515,
input WL516,
input WL517,
input WL518,
input WL519,
input WL520,
input WL521,
input WL522,
input WL523,
input WL524,
input WL525,
input WL526,
input WL527,
input WL528,
input WL529,
input WL530,
input WL531,
input WL532,
input WL533,
input WL534,
input WL535,
input WL536,
input WL537,
input WL538,
input WL539,
input WL540,
input WL541,
input WL542,
input WL543,
input WL544,
input WL545,
input WL546,
input WL547,
input WL548,
input WL549,
input WL550,
input WL551,
input WL552,
input WL553,
input WL554,
input WL555,
input WL556,
input WL557,
input WL558,
input WL559,
input WL560,
input WL561,
input WL562,
input WL563,
input WL564,
input WL565,
input WL566,
input WL567,
input WL568,
input WL569,
input WL570,
input WL571,
input WL572,
input WL573,
input WL574,
input WL575,
input WL576,
input WL577,
input WL578,
input WL579,
input WL580,
input WL581,
input WL582,
input WL583,
input WL584,
input WL585,
input WL586,
input WL587,
input WL588,
input WL589,
input WL590,
input WL591,
input WL592,
input WL593,
input WL594,
input WL595,
input WL596,
input WL597,
input WL598,
input WL599,
input WL600,
input WL601,
input WL602,
input WL603,
input WL604,
input WL605,
input WL606,
input WL607,
input WL608,
input WL609,
input WL610,
input WL611,
input WL612,
input WL613,
input WL614,
input WL615,
input WL616,
input WL617,
input WL618,
input WL619,
input WL620,
input WL621,
input WL622,
input WL623,
input WL624,
input WL625,
input WL626,
input WL627,
input WL628,
input WL629,
input WL630,
input WL631,
input WL632,
input WL633,
input WL634,
input WL635,
input WL636,
input WL637,
input WL638,
input WL639,
input WL640,
input WL641,
input WL642,
input WL643,
input WL644,
input WL645,
input WL646,
input WL647,
input WL648,
input WL649,
input WL650,
input WL651,
input WL652,
input WL653,
input WL654,
input WL655,
input WL656,
input WL657,
input WL658,
input WL659,
input WL660,
input WL661,
input WL662,
input WL663,
input WL664,
input WL665,
input WL666,
input WL667,
input WL668,
input WL669,
input WL670,
input WL671,
input WL672,
input WL673,
input WL674,
input WL675,
input WL676,
input WL677,
input WL678,
input WL679,
input WL680,
input WL681,
input WL682,
input WL683,
input WL684,
input WL685,
input WL686,
input WL687,
input WL688,
input WL689,
input WL690,
input WL691,
input WL692,
input WL693,
input WL694,
input WL695,
input WL696,
input WL697,
input WL698,
input WL699,
input WL700,
input WL701,
input WL702,
input WL703,
input WL704,
input WL705,
input WL706,
input WL707,
input WL708,
input WL709,
input WL710,
input WL711,
input WL712,
input WL713,
input WL714,
input WL715,
input WL716,
input WL717,
input WL718,
input WL719,
input WL720,
input WL721,
input WL722,
input WL723,
input WL724,
input WL725,
input WL726,
input WL727,
input WL728,
input WL729,
input WL730,
input WL731,
input WL732,
input WL733,
input WL734,
input WL735,
input WL736,
input WL737,
input WL738,
input WL739,
input WL740,
input WL741,
input WL742,
input WL743,
input WL744,
input WL745,
input WL746,
input WL747,
input WL748,
input WL749,
input WL750,
input WL751,
input WL752,
input WL753,
input WL754,
input WL755,
input WL756,
input WL757,
input WL758,
input WL759,
input WL760,
input WL761,
input WL762,
input WL763,
input WL764,
input WL765,
input WL766,
input WL767,
input WL768,
input WL769,
input WL770,
input WL771,
input WL772,
input WL773,
input WL774,
input WL775,
input WL776,
input WL777,
input WL778,
input WL779,
input WL780,
input WL781,
input WL782,
input WL783,
input WL784,
input WL785,
input WL786,
input WL787,
input WL788,
input WL789,
input WL790,
input WL791,
input WL792,
input WL793,
input WL794,
input WL795,
input WL796,
input WL797,
input WL798,
input WL799,
input WL800,
input WL801,
input WL802,
input WL803,
input WL804,
input WL805,
input WL806,
input WL807,
input WL808,
input WL809,
input WL810,
input WL811,
input WL812,
input WL813,
input WL814,
input WL815,
input WL816,
input WL817,
input WL818,
input WL819,
input WL820,
input WL821,
input WL822,
input WL823,
input WL824,
input WL825,
input WL826,
input WL827,
input WL828,
input WL829,
input WL830,
input WL831,
input WL832,
input WL833,
input WL834,
input WL835,
input WL836,
input WL837,
input WL838,
input WL839,
input WL840,
input WL841,
input WL842,
input WL843,
input WL844,
input WL845,
input WL846,
input WL847,
input WL848,
input WL849,
input WL850,
input WL851,
input WL852,
input WL853,
input WL854,
input WL855,
input WL856,
input WL857,
input WL858,
input WL859,
input WL860,
input WL861,
input WL862,
input WL863,
input WL864,
input WL865,
input WL866,
input WL867,
input WL868,
input WL869,
input WL870,
input WL871,
input WL872,
input WL873,
input WL874,
input WL875,
input WL876,
input WL877,
input WL878,
input WL879,
input WL880,
input WL881,
input WL882,
input WL883,
input WL884,
input WL885,
input WL886,
input WL887,
input WL888,
input WL889,
input WL890,
input WL891,
input WL892,
input WL893,
input WL894,
input WL895,
input WL896,
input WL897,
input WL898,
input WL899,
input WL900,
input WL901,
input WL902,
input WL903,
input WL904,
input WL905,
input WL906,
input WL907,
input WL908,
input WL909,
input WL910,
input WL911,
input WL912,
input WL913,
input WL914,
input WL915,
input WL916,
input WL917,
input WL918,
input WL919,
input WL920,
input WL921,
input WL922,
input WL923,
input WL924,
input WL925,
input WL926,
input WL927,
input WL928,
input WL929,
input WL930,
input WL931,
input WL932,
input WL933,
input WL934,
input WL935,
input WL936,
input WL937,
input WL938,
input WL939,
input WL940,
input WL941,
input WL942,
input WL943,
input WL944,
input WL945,
input WL946,
input WL947,
input WL948,
input WL949,
input WL950,
input WL951,
input WL952,
input WL953,
input WL954,
input WL955,
input WL956,
input WL957,
input WL958,
input WL959,
input WL960,
input WL961,
input WL962,
input WL963,
input WL964,
input WL965,
input WL966,
input WL967,
input WL968,
input WL969,
input WL970,
input WL971,
input WL972,
input WL973,
input WL974,
input WL975,
input WL976,
input WL977,
input WL978,
input WL979,
input WL980,
input WL981,
input WL982,
input WL983,
input WL984,
input WL985,
input WL986,
input WL987,
input WL988,
input WL989,
input WL990,
input WL991,
input WL992,
input WL993,
input WL994,
input WL995,
input WL996,
input WL997,
input WL998,
input WL999,
input WL1000,
input WL1001,
input WL1002,
input WL1003,
input WL1004,
input WL1005,
input WL1006,
input WL1007,
input WL1008,
input WL1009,
input WL1010,
input WL1011,
input WL1012,
input WL1013,
input WL1014,
input WL1015,
input WL1016,
input WL1017,
input WL1018,
input WL1019,
input WL1020,
input WL1021,
input WL1022,
input WL1023

   
);
endmodule
`default_nettype wire
