// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

module data_in_decoder (
		input [7:0] data_in,
                input [1:0] sel,
                output reg [31:0] data_out
);

always @(*) begin
   case (sel)
      2'b00: data_out[7:0] = data_in;
      2'b01: data_out[15:8] = data_in;
      2'b10: data_out[23:16] = data_in;
      2'b11: data_out[32:24] = data_in;
   endcase
end

endmodule
