VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj_IMPACT_HEAD
  CLASS BLOCK ;
  FOREIGN user_proj_IMPACT_HEAD ;
  ORIGIN 0.000 0.000 ;
  SIZE 800.000 BY 760.000 ;
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 4.000 40.080 ;
    END
  END C
  PIN East[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 107.480 4.000 108.080 ;
    END
  END East[0]
  PIN East[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 175.480 4.000 176.080 ;
    END
  END East[1]
  PIN East[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 243.480 4.000 244.080 ;
    END
  END East[2]
  PIN East[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 311.480 4.000 312.080 ;
    END
  END East[3]
  PIN East[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 379.480 4.000 380.080 ;
    END
  END East[4]
  PIN East[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 447.480 4.000 448.080 ;
    END
  END East[5]
  PIN East[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 515.480 4.000 516.080 ;
    END
  END East[6]
  PIN East[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 583.480 4.000 584.080 ;
    END
  END East[7]
  PIN East[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 651.480 4.000 652.080 ;
    END
  END East[8]
  PIN East[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 719.480 4.000 720.080 ;
    END
  END East[9]
  PIN PO[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.383400 ;
    PORT
      LAYER met3 ;
        RECT 796.000 42.200 800.000 42.800 ;
    END
  END PO[0]
  PIN PO[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.383400 ;
    PORT
      LAYER met3 ;
        RECT 796.000 126.520 800.000 127.120 ;
    END
  END PO[1]
  PIN PO[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.383400 ;
    PORT
      LAYER met3 ;
        RECT 796.000 210.840 800.000 211.440 ;
    END
  END PO[2]
  PIN PO[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.383400 ;
    PORT
      LAYER met3 ;
        RECT 796.000 295.160 800.000 295.760 ;
    END
  END PO[3]
  PIN PO[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.383400 ;
    PORT
      LAYER met3 ;
        RECT 796.000 379.480 800.000 380.080 ;
    END
  END PO[4]
  PIN PO[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.383400 ;
    PORT
      LAYER met3 ;
        RECT 796.000 463.800 800.000 464.400 ;
    END
  END PO[5]
  PIN PO[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.383400 ;
    PORT
      LAYER met3 ;
        RECT 796.000 548.120 800.000 548.720 ;
    END
  END PO[6]
  PIN PO[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.383400 ;
    PORT
      LAYER met3 ;
        RECT 796.000 632.440 800.000 633.040 ;
    END
  END PO[7]
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 36.430 0.000 36.710 4.000 ;
    END
  END SI
  PIN WL_Bank01[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.383400 ;
    PORT
      LAYER met2 ;
        RECT 109.110 0.000 109.390 4.000 ;
    END
  END WL_Bank01[0]
  PIN WL_Bank01[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.383400 ;
    PORT
      LAYER met2 ;
        RECT 181.790 0.000 182.070 4.000 ;
    END
  END WL_Bank01[1]
  PIN WL_Bank01[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.383400 ;
    PORT
      LAYER met2 ;
        RECT 254.470 0.000 254.750 4.000 ;
    END
  END WL_Bank01[2]
  PIN WL_Bank01[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.383400 ;
    PORT
      LAYER met2 ;
        RECT 327.150 0.000 327.430 4.000 ;
    END
  END WL_Bank01[3]
  PIN WL_Bank01[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.383400 ;
    PORT
      LAYER met2 ;
        RECT 399.830 0.000 400.110 4.000 ;
    END
  END WL_Bank01[4]
  PIN WL_Bank01[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.383400 ;
    PORT
      LAYER met2 ;
        RECT 472.510 0.000 472.790 4.000 ;
    END
  END WL_Bank01[5]
  PIN WL_Bank01[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.383400 ;
    PORT
      LAYER met2 ;
        RECT 545.190 0.000 545.470 4.000 ;
    END
  END WL_Bank01[6]
  PIN WL_Bank01[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.383400 ;
    PORT
      LAYER met2 ;
        RECT 617.870 0.000 618.150 4.000 ;
    END
  END WL_Bank01[7]
  PIN WL_Bank01[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.383400 ;
    PORT
      LAYER met2 ;
        RECT 690.550 0.000 690.830 4.000 ;
    END
  END WL_Bank01[8]
  PIN WL_Bank01[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.383400 ;
    PORT
      LAYER met2 ;
        RECT 763.230 0.000 763.510 4.000 ;
    END
  END WL_Bank01[9]
  PIN test
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 716.760 800.000 717.360 ;
    END
  END test
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 748.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 748.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 748.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 748.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 748.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 748.240 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 748.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 748.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 748.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 748.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 748.240 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 794.420 748.085 ;
      LAYER met1 ;
        RECT 4.670 10.240 794.420 748.240 ;
      LAYER met2 ;
        RECT 4.690 4.280 792.950 748.185 ;
        RECT 4.690 4.000 36.150 4.280 ;
        RECT 36.990 4.000 108.830 4.280 ;
        RECT 109.670 4.000 181.510 4.280 ;
        RECT 182.350 4.000 254.190 4.280 ;
        RECT 255.030 4.000 326.870 4.280 ;
        RECT 327.710 4.000 399.550 4.280 ;
        RECT 400.390 4.000 472.230 4.280 ;
        RECT 473.070 4.000 544.910 4.280 ;
        RECT 545.750 4.000 617.590 4.280 ;
        RECT 618.430 4.000 690.270 4.280 ;
        RECT 691.110 4.000 762.950 4.280 ;
        RECT 763.790 4.000 792.950 4.280 ;
      LAYER met3 ;
        RECT 3.990 720.480 796.000 748.165 ;
        RECT 4.400 719.080 796.000 720.480 ;
        RECT 3.990 717.760 796.000 719.080 ;
        RECT 3.990 716.360 795.600 717.760 ;
        RECT 3.990 652.480 796.000 716.360 ;
        RECT 4.400 651.080 796.000 652.480 ;
        RECT 3.990 633.440 796.000 651.080 ;
        RECT 3.990 632.040 795.600 633.440 ;
        RECT 3.990 584.480 796.000 632.040 ;
        RECT 4.400 583.080 796.000 584.480 ;
        RECT 3.990 549.120 796.000 583.080 ;
        RECT 3.990 547.720 795.600 549.120 ;
        RECT 3.990 516.480 796.000 547.720 ;
        RECT 4.400 515.080 796.000 516.480 ;
        RECT 3.990 464.800 796.000 515.080 ;
        RECT 3.990 463.400 795.600 464.800 ;
        RECT 3.990 448.480 796.000 463.400 ;
        RECT 4.400 447.080 796.000 448.480 ;
        RECT 3.990 380.480 796.000 447.080 ;
        RECT 4.400 379.080 795.600 380.480 ;
        RECT 3.990 312.480 796.000 379.080 ;
        RECT 4.400 311.080 796.000 312.480 ;
        RECT 3.990 296.160 796.000 311.080 ;
        RECT 3.990 294.760 795.600 296.160 ;
        RECT 3.990 244.480 796.000 294.760 ;
        RECT 4.400 243.080 796.000 244.480 ;
        RECT 3.990 211.840 796.000 243.080 ;
        RECT 3.990 210.440 795.600 211.840 ;
        RECT 3.990 176.480 796.000 210.440 ;
        RECT 4.400 175.080 796.000 176.480 ;
        RECT 3.990 127.520 796.000 175.080 ;
        RECT 3.990 126.120 795.600 127.520 ;
        RECT 3.990 108.480 796.000 126.120 ;
        RECT 4.400 107.080 796.000 108.480 ;
        RECT 3.990 43.200 796.000 107.080 ;
        RECT 3.990 41.800 795.600 43.200 ;
        RECT 3.990 40.480 796.000 41.800 ;
        RECT 4.400 39.080 796.000 40.480 ;
        RECT 3.990 10.715 796.000 39.080 ;
  END
END user_proj_IMPACT_HEAD
END LIBRARY

