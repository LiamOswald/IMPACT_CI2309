VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj_IMPACT_HEAD
  CLASS BLOCK ;
  FOREIGN user_proj_IMPACT_HEAD ;
  ORIGIN 0.000 0.000 ;
  SIZE 2400.000 BY 3000.000 ;
  PIN Bank_Select[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 375.400 4.000 376.000 ;
    END
  END Bank_Select[0]
  PIN Bank_Select[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1124.760 4.000 1125.360 ;
    END
  END Bank_Select[1]
  PIN Byte_Select[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1874.120 4.000 1874.720 ;
    END
  END Byte_Select[0]
  PIN Byte_Select[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2623.480 4.000 2624.080 ;
    END
  END Byte_Select[1]
  PIN Data_In[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 75.070 0.000 75.350 4.000 ;
    END
  END Data_In[0]
  PIN Data_In[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 225.030 0.000 225.310 4.000 ;
    END
  END Data_In[1]
  PIN Data_In[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 374.990 0.000 375.270 4.000 ;
    END
  END Data_In[2]
  PIN Data_In[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 524.950 0.000 525.230 4.000 ;
    END
  END Data_In[3]
  PIN Data_In[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 674.910 0.000 675.190 4.000 ;
    END
  END Data_In[4]
  PIN Data_In[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 824.870 0.000 825.150 4.000 ;
    END
  END Data_In[5]
  PIN Data_In[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 974.830 0.000 975.110 4.000 ;
    END
  END Data_In[6]
  PIN Data_In[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 1124.790 0.000 1125.070 4.000 ;
    END
  END Data_In[7]
  PIN Data_Out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.383400 ;
    PORT
      LAYER met2 ;
        RECT 1274.750 0.000 1275.030 4.000 ;
    END
  END Data_Out[0]
  PIN Data_Out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.383400 ;
    PORT
      LAYER met2 ;
        RECT 1424.710 0.000 1424.990 4.000 ;
    END
  END Data_Out[1]
  PIN Data_Out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.383400 ;
    PORT
      LAYER met2 ;
        RECT 1574.670 0.000 1574.950 4.000 ;
    END
  END Data_Out[2]
  PIN Data_Out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.383400 ;
    PORT
      LAYER met2 ;
        RECT 1724.630 0.000 1724.910 4.000 ;
    END
  END Data_Out[3]
  PIN Data_Out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.383400 ;
    PORT
      LAYER met2 ;
        RECT 1874.590 0.000 1874.870 4.000 ;
    END
  END Data_Out[4]
  PIN Data_Out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.383400 ;
    PORT
      LAYER met2 ;
        RECT 2024.550 0.000 2024.830 4.000 ;
    END
  END Data_Out[5]
  PIN Data_Out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.383400 ;
    PORT
      LAYER met2 ;
        RECT 2174.510 0.000 2174.790 4.000 ;
    END
  END Data_Out[6]
  PIN Data_Out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.383400 ;
    PORT
      LAYER met2 ;
        RECT 2324.470 0.000 2324.750 4.000 ;
    END
  END Data_Out[7]
  PIN PreCharge
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 201.570 2996.000 201.850 3000.000 ;
    END
  END PreCharge
  PIN ReadEnable
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 87.490 2996.000 87.770 3000.000 ;
    END
  END ReadEnable
  PIN Word_Select[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2396.000 152.360 2400.000 152.960 ;
    END
  END Word_Select[0]
  PIN Word_Select[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2396.000 451.560 2400.000 452.160 ;
    END
  END Word_Select[1]
  PIN Word_Select[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 2396.000 750.760 2400.000 751.360 ;
    END
  END Word_Select[2]
  PIN Word_Select[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 2396.000 1049.960 2400.000 1050.560 ;
    END
  END Word_Select[3]
  PIN Word_Select[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2396.000 1349.160 2400.000 1349.760 ;
    END
  END Word_Select[4]
  PIN Word_Select[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 2396.000 1648.360 2400.000 1648.960 ;
    END
  END Word_Select[5]
  PIN Word_Select[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 2396.000 1947.560 2400.000 1948.160 ;
    END
  END Word_Select[6]
  PIN Word_Select[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2396.000 2246.760 2400.000 2247.360 ;
    END
  END Word_Select[7]
  PIN Word_Select[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2396.000 2545.960 2400.000 2546.560 ;
    END
  END Word_Select[8]
  PIN Word_Select[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met3 ;
        RECT 2396.000 2845.160 2400.000 2845.760 ;
    END
  END Word_Select[9]
  PIN WriteEnable
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 30.450 2996.000 30.730 3000.000 ;
    END
  END WriteEnable
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 144.530 2996.000 144.810 3000.000 ;
    END
  END clk
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.610 2996.000 258.890 3000.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 829.010 2996.000 829.290 3000.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 886.050 2996.000 886.330 3000.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 943.090 2996.000 943.370 3000.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1000.130 2996.000 1000.410 3000.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1057.170 2996.000 1057.450 3000.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1114.210 2996.000 1114.490 3000.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1171.250 2996.000 1171.530 3000.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1228.290 2996.000 1228.570 3000.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1285.330 2996.000 1285.610 3000.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1342.370 2996.000 1342.650 3000.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 2996.000 315.930 3000.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1399.410 2996.000 1399.690 3000.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1456.450 2996.000 1456.730 3000.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1513.490 2996.000 1513.770 3000.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1570.530 2996.000 1570.810 3000.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1627.570 2996.000 1627.850 3000.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1684.610 2996.000 1684.890 3000.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1741.650 2996.000 1741.930 3000.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1798.690 2996.000 1798.970 3000.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1855.730 2996.000 1856.010 3000.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1912.770 2996.000 1913.050 3000.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.690 2996.000 372.970 3000.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1969.810 2996.000 1970.090 3000.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2026.850 2996.000 2027.130 3000.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2083.890 2996.000 2084.170 3000.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2140.930 2996.000 2141.210 3000.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2197.970 2996.000 2198.250 3000.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2255.010 2996.000 2255.290 3000.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2312.050 2996.000 2312.330 3000.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2369.090 2996.000 2369.370 3000.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 429.730 2996.000 430.010 3000.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.770 2996.000 487.050 3000.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.810 2996.000 544.090 3000.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 600.850 2996.000 601.130 3000.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 657.890 2996.000 658.170 3000.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.930 2996.000 715.210 3000.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.970 2996.000 772.250 3000.000 ;
    END
  END io_oeb[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 451.415 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 2697.225 944.240 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 451.415 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 2697.225 1097.840 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 451.415 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 2697.225 1251.440 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 451.415 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 2697.225 1405.040 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.040 10.640 1558.640 451.415 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.040 2697.225 1558.640 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1710.640 10.640 1712.240 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1864.240 10.640 1865.840 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2017.840 10.640 2019.440 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2171.440 10.640 2173.040 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2325.040 10.640 2326.640 2986.800 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 451.415 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 2697.225 867.440 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 451.415 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 2697.225 1021.040 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 451.415 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 2697.225 1174.640 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 451.415 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 2697.225 1328.240 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 451.415 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 2697.225 1481.840 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1633.840 10.640 1635.440 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1787.440 10.640 1789.040 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 1941.040 10.640 1942.640 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2094.640 10.640 2096.240 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2248.240 10.640 2249.840 2986.800 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2394.300 2986.645 ;
      LAYER met1 ;
        RECT 4.670 10.640 2394.300 2986.800 ;
      LAYER met2 ;
        RECT 4.690 2995.720 30.170 2996.490 ;
        RECT 31.010 2995.720 87.210 2996.490 ;
        RECT 88.050 2995.720 144.250 2996.490 ;
        RECT 145.090 2995.720 201.290 2996.490 ;
        RECT 202.130 2995.720 258.330 2996.490 ;
        RECT 259.170 2995.720 315.370 2996.490 ;
        RECT 316.210 2995.720 372.410 2996.490 ;
        RECT 373.250 2995.720 429.450 2996.490 ;
        RECT 430.290 2995.720 486.490 2996.490 ;
        RECT 487.330 2995.720 543.530 2996.490 ;
        RECT 544.370 2995.720 600.570 2996.490 ;
        RECT 601.410 2995.720 657.610 2996.490 ;
        RECT 658.450 2995.720 714.650 2996.490 ;
        RECT 715.490 2995.720 771.690 2996.490 ;
        RECT 772.530 2995.720 828.730 2996.490 ;
        RECT 829.570 2995.720 885.770 2996.490 ;
        RECT 886.610 2995.720 942.810 2996.490 ;
        RECT 943.650 2995.720 999.850 2996.490 ;
        RECT 1000.690 2995.720 1056.890 2996.490 ;
        RECT 1057.730 2995.720 1113.930 2996.490 ;
        RECT 1114.770 2995.720 1170.970 2996.490 ;
        RECT 1171.810 2995.720 1228.010 2996.490 ;
        RECT 1228.850 2995.720 1285.050 2996.490 ;
        RECT 1285.890 2995.720 1342.090 2996.490 ;
        RECT 1342.930 2995.720 1399.130 2996.490 ;
        RECT 1399.970 2995.720 1456.170 2996.490 ;
        RECT 1457.010 2995.720 1513.210 2996.490 ;
        RECT 1514.050 2995.720 1570.250 2996.490 ;
        RECT 1571.090 2995.720 1627.290 2996.490 ;
        RECT 1628.130 2995.720 1684.330 2996.490 ;
        RECT 1685.170 2995.720 1741.370 2996.490 ;
        RECT 1742.210 2995.720 1798.410 2996.490 ;
        RECT 1799.250 2995.720 1855.450 2996.490 ;
        RECT 1856.290 2995.720 1912.490 2996.490 ;
        RECT 1913.330 2995.720 1969.530 2996.490 ;
        RECT 1970.370 2995.720 2026.570 2996.490 ;
        RECT 2027.410 2995.720 2083.610 2996.490 ;
        RECT 2084.450 2995.720 2140.650 2996.490 ;
        RECT 2141.490 2995.720 2197.690 2996.490 ;
        RECT 2198.530 2995.720 2254.730 2996.490 ;
        RECT 2255.570 2995.720 2311.770 2996.490 ;
        RECT 2312.610 2995.720 2368.810 2996.490 ;
        RECT 2369.650 2995.720 2393.290 2996.490 ;
        RECT 4.690 4.280 2393.290 2995.720 ;
        RECT 4.690 3.670 74.790 4.280 ;
        RECT 75.630 3.670 224.750 4.280 ;
        RECT 225.590 3.670 374.710 4.280 ;
        RECT 375.550 3.670 524.670 4.280 ;
        RECT 525.510 3.670 674.630 4.280 ;
        RECT 675.470 3.670 824.590 4.280 ;
        RECT 825.430 3.670 974.550 4.280 ;
        RECT 975.390 3.670 1124.510 4.280 ;
        RECT 1125.350 3.670 1274.470 4.280 ;
        RECT 1275.310 3.670 1424.430 4.280 ;
        RECT 1425.270 3.670 1574.390 4.280 ;
        RECT 1575.230 3.670 1724.350 4.280 ;
        RECT 1725.190 3.670 1874.310 4.280 ;
        RECT 1875.150 3.670 2024.270 4.280 ;
        RECT 2025.110 3.670 2174.230 4.280 ;
        RECT 2175.070 3.670 2324.190 4.280 ;
        RECT 2325.030 3.670 2393.290 4.280 ;
      LAYER met3 ;
        RECT 4.000 2846.160 2396.000 2986.725 ;
        RECT 4.000 2844.760 2395.600 2846.160 ;
        RECT 4.000 2624.480 2396.000 2844.760 ;
        RECT 4.400 2623.080 2396.000 2624.480 ;
        RECT 4.000 2546.960 2396.000 2623.080 ;
        RECT 4.000 2545.560 2395.600 2546.960 ;
        RECT 4.000 2247.760 2396.000 2545.560 ;
        RECT 4.000 2246.360 2395.600 2247.760 ;
        RECT 4.000 1948.560 2396.000 2246.360 ;
        RECT 4.000 1947.160 2395.600 1948.560 ;
        RECT 4.000 1875.120 2396.000 1947.160 ;
        RECT 4.400 1873.720 2396.000 1875.120 ;
        RECT 4.000 1649.360 2396.000 1873.720 ;
        RECT 4.000 1647.960 2395.600 1649.360 ;
        RECT 4.000 1350.160 2396.000 1647.960 ;
        RECT 4.000 1348.760 2395.600 1350.160 ;
        RECT 4.000 1125.760 2396.000 1348.760 ;
        RECT 4.400 1124.360 2396.000 1125.760 ;
        RECT 4.000 1050.960 2396.000 1124.360 ;
        RECT 4.000 1049.560 2395.600 1050.960 ;
        RECT 4.000 751.760 2396.000 1049.560 ;
        RECT 4.000 750.360 2395.600 751.760 ;
        RECT 4.000 452.560 2396.000 750.360 ;
        RECT 4.000 451.160 2395.600 452.560 ;
        RECT 4.000 376.400 2396.000 451.160 ;
        RECT 4.400 375.000 2396.000 376.400 ;
        RECT 4.000 153.360 2396.000 375.000 ;
        RECT 4.000 151.960 2395.600 153.360 ;
        RECT 4.000 10.715 2396.000 151.960 ;
      LAYER met4 ;
        RECT 751.015 11.735 788.640 2723.905 ;
        RECT 791.040 2696.825 865.440 2723.905 ;
        RECT 867.840 2696.825 942.240 2723.905 ;
        RECT 944.640 2696.825 1019.040 2723.905 ;
        RECT 1021.440 2696.825 1095.840 2723.905 ;
        RECT 1098.240 2696.825 1172.640 2723.905 ;
        RECT 1175.040 2696.825 1249.440 2723.905 ;
        RECT 1251.840 2696.825 1326.240 2723.905 ;
        RECT 1328.640 2696.825 1403.040 2723.905 ;
        RECT 1405.440 2696.825 1479.840 2723.905 ;
        RECT 1482.240 2696.825 1556.640 2723.905 ;
        RECT 1559.040 2696.825 1633.440 2723.905 ;
        RECT 791.040 451.815 1633.440 2696.825 ;
        RECT 791.040 11.735 865.440 451.815 ;
        RECT 867.840 11.735 942.240 451.815 ;
        RECT 944.640 11.735 1019.040 451.815 ;
        RECT 1021.440 11.735 1095.840 451.815 ;
        RECT 1098.240 11.735 1172.640 451.815 ;
        RECT 1175.040 11.735 1249.440 451.815 ;
        RECT 1251.840 11.735 1326.240 451.815 ;
        RECT 1328.640 11.735 1403.040 451.815 ;
        RECT 1405.440 11.735 1479.840 451.815 ;
        RECT 1482.240 11.735 1556.640 451.815 ;
        RECT 1559.040 11.735 1633.440 451.815 ;
        RECT 1635.840 11.735 1657.545 2723.905 ;
  END
END user_proj_IMPACT_HEAD
END LIBRARY

