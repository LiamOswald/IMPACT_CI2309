
/*
// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0
 *-------------------------------------------------------------
 *
 * user_proj_IMPACT_Head
 * 
 * This head was built by LiamOswald for the University of South Alabama's SRAM research into various SRAM banks
 * If Liam isn't lazy, he will update this comment with real information at a later date... don't bet on it. 
 * Email him: wdo1621@jagmail.southalabama.edu
 *
 *-------------------------------------------------------------
 */
 `default_nettype none
`include "user_defines.v"

module user_proj_IMPACT_HEAD (

`ifdef USE_POWER_PINS
    inout vccd1,	// User area 1 1.8V supply
    inout vssd1,	// User area 1 digital ground
`endif

output [37:0] io_oeb,
    // IRQ
output wire [2:0] user_irq,
input wire [7:0] Data_In,				//SRAM byte input		GPIO pins 0-7
output wire [7:0] Data_Out, 				//SRAM byte output		GPIO pins 8-15
input wire [9:0] Word_Select,				/////////////////////////////////////changed 9 to 4///////////////////////////
//input wire [1:0] Bank_Select, 				//Select SRAM Bank		GPIO pins 26 & 27
input wire [1:0] Byte_Select, 				//Select Byte from Word		GPIO pins 28 & 29
input wire WriteEnable,					//SRAM Write Enable signal	GPIO pin 30
input wire ReadEnable,
input wire WL_enable,					//SRAM Read Enable Signal	GPIO pin 31
input wire PreCharge,
input clk					//PreCharge	GPIO pin 32
);

assign io_oeb = 38'b11111111_00000000_1111111111_11_11_1_1_0_11_10_1;
assign user_irq = 3'b000;	// Unused

wire [31:0] SRAM_In;
			
wire [1023:0] WL;		///////////////////////////changed 1023 to 31 if 32 by 32 sram
wire [31:0] SRAM_Out;




//################################################
//Creates the Four Word Decoders Instences for the Four Memory Banks
//################################################

// BANK 01 WORDLINE Decoder
BankWordDecoder wordDecoder_Bank01 (
	.clk(clk),
	.sel(Word_Select),
	.WL_enable(WL_enable),
	.address(WL)
);

//DATA OUT MUX! this mux takes 4 32bit values from the 4 memory banks, and mux's the output down to a single byte ready for the output pins
OneBankMux Data_out_Mux(
		.clk(clk),
		.read_enable(ReadEnable),
		.Bank01_Reading(SRAM_Out),	
		.byte_sel(Byte_Select),
                .data_out(Data_Out)
);

data_in_decoder DataIn_Decoder(
	.clk(clk),
	.write_enable(WriteEnable),
	.data_in(Data_In),
	.sel(Byte_Select),
	.data_out(SRAM_In)
);


//BANKBANKBANKBANKBANKBANKBANKBANKBANKBANKBANKBANKBANKBANKBANKBANKBANKBANKBANKBANKBANKBANKBANKBANKBANKBANKBANKBANK
//BANKBANKBANKBANKBANKBA     bank                                       NKBANKBANKBANKBANKBANKBANKBANKBANKBANKBANK
//BANKBANKBANKBANKBANKBANKBANKBANKBANKBANKBANKBANKBANKBANKBANKBANKBANKBANKBANKBANKBANKBANKBANKBANKBANKBANKBANKBANK

//Bank01 SRAM Block
full_sram bank01(      
	
	`ifdef USE_POWER_PINS
    		.vccd1(vccd1),	// User area 1 1.8V supply
    		.vssd1(vssd1),	// User area 1 digital ground
	`endif
	
.PRE(PreCharge),
.readen(ReadEnable),
.writeen(WriteEnable),

.DataIn0(SRAM_In [0]),
.DataIn1(SRAM_In [1]),
.DataIn2(SRAM_In [2]),
.DataIn3(SRAM_In [3]),
.DataIn4(SRAM_In [4]),
.DataIn5(SRAM_In [5]),
.DataIn6(SRAM_In [6]),
.DataIn7(SRAM_In [7]),
.DataIn8(SRAM_In [8]),
.DataIn9(SRAM_In [9]),
.DataIn10(SRAM_In [10]),
.DataIn11(SRAM_In [11]),
.DataIn12(SRAM_In [12]),
.DataIn13(SRAM_In [13]),
.DataIn14(SRAM_In [14]),
.DataIn15(SRAM_In [15]),
.DataIn16(SRAM_In [16]),
.DataIn17(SRAM_In [17]),
.DataIn18(SRAM_In [18]),
.DataIn19(SRAM_In [19]),
.DataIn20(SRAM_In [20]),
.DataIn21(SRAM_In [21]),
.DataIn22(SRAM_In [22]),
.DataIn23(SRAM_In [23]),
.DataIn24(SRAM_In [24]),
.DataIn25(SRAM_In [25]),
.DataIn26(SRAM_In [26]),
.DataIn27(SRAM_In [27]),
.DataIn28(SRAM_In [28]),
.DataIn29(SRAM_In [29]),
.DataIn30(SRAM_In [30]),
.DataIn31(SRAM_In [31]),


.DataOut0(SRAM_Out [0]),
.DataOut1(SRAM_Out [1]),
.DataOut2(SRAM_Out [2]),
.DataOut3(SRAM_Out [3]),
.DataOut4(SRAM_Out [4]),
.DataOut5(SRAM_Out [5]),
.DataOut6(SRAM_Out [6]),
.DataOut7(SRAM_Out [7]),
.DataOut8(SRAM_Out [8]),
.DataOut9(SRAM_Out [9]),
.DataOut10(SRAM_Out [10]),
.DataOut11(SRAM_Out [11]),
.DataOut12(SRAM_Out [12]),
.DataOut13(SRAM_Out [13]),
.DataOut14(SRAM_Out [14]),
.DataOut15(SRAM_Out [15]),
.DataOut16(SRAM_Out [16]),
.DataOut17(SRAM_Out [17]),
.DataOut18(SRAM_Out [18]),
.DataOut19(SRAM_Out [19]),
.DataOut20(SRAM_Out [20]),
.DataOut21(SRAM_Out [21]),
.DataOut22(SRAM_Out [22]),
.DataOut23(SRAM_Out [23]),
.DataOut24(SRAM_Out [24]),
.DataOut25(SRAM_Out [25]),
.DataOut26(SRAM_Out [26]),
.DataOut27(SRAM_Out [27]),
.DataOut28(SRAM_Out [28]),
.DataOut29(SRAM_Out [29]),
.DataOut30(SRAM_Out [30]),
.DataOut31(SRAM_Out [31]),


.WL0(WL [0]),
.WL1(WL [1]),
.WL2(WL [2]),
.WL3(WL [3]),
.WL4(WL [4]),
.WL5(WL [5]),
.WL6(WL [6]),
.WL7(WL [7]),
.WL8(WL [8]),
.WL9(WL [9]),
.WL10(WL [10]),
.WL11(WL [11]),
.WL12(WL [12]),
.WL13(WL [13]),
.WL14(WL [14]),
.WL15(WL [15]),
.WL16(WL [16]),
.WL17(WL [17]),
.WL18(WL [18]),
.WL19(WL [19]),
.WL20(WL [20]),
.WL21(WL [21]),
.WL22(WL [22]),
.WL23(WL [23]),
.WL24(WL [24]),
.WL25(WL [25]),
.WL26(WL [26]),
.WL27(WL [27]),
.WL28(WL [28]),
.WL29(WL [29]),
.WL30(WL [30]),
.WL31(WL [31]),
.WL32(WL [32]),
.WL33(WL [33]),
.WL34(WL [34]),
.WL35(WL [35]),
.WL36(WL [36]),
.WL37(WL [37]),
.WL38(WL [38]),
.WL39(WL [39]),
.WL40(WL [40]),
.WL41(WL [41]),
.WL42(WL [42]),
.WL43(WL [43]),
.WL44(WL [44]),
.WL45(WL [45]),
.WL46(WL [46]),
.WL47(WL [47]),
.WL48(WL [48]),
.WL49(WL [49]),
.WL50(WL [50]),
.WL51(WL [51]),
.WL52(WL [52]),
.WL53(WL [53]),
.WL54(WL [54]),
.WL55(WL [55]),
.WL56(WL [56]),
.WL57(WL [57]),
.WL58(WL [58]),
.WL59(WL [59]),
.WL60(WL [60]),
.WL61(WL [61]),
.WL62(WL [62]),
.WL63(WL [63]),
.WL64(WL [64]),
.WL65(WL [65]),
.WL66(WL [66]),
.WL67(WL [67]),
.WL68(WL [68]),
.WL69(WL [69]),
.WL70(WL [70]),
.WL71(WL [71]),
.WL72(WL [72]),
.WL73(WL [73]),
.WL74(WL [74]),
.WL75(WL [75]),
.WL76(WL [76]),
.WL77(WL [77]),
.WL78(WL [78]),
.WL79(WL [79]),
.WL80(WL [80]),
.WL81(WL [81]),
.WL82(WL [82]),
.WL83(WL [83]),
.WL84(WL [84]),
.WL85(WL [85]),
.WL86(WL [86]),
.WL87(WL [87]),
.WL88(WL [88]),
.WL89(WL [89]),
.WL90(WL [90]),
.WL91(WL [91]),
.WL92(WL [92]),
.WL93(WL [93]),
.WL94(WL [94]),
.WL95(WL [95]),
.WL96(WL [96]),
.WL97(WL [97]),
.WL98(WL [98]),
.WL99(WL [99]),
.WL100(WL [100]),
.WL101(WL [101]),
.WL102(WL [102]),
.WL103(WL [103]),
.WL104(WL [104]),
.WL105(WL [105]),
.WL106(WL [106]),
.WL107(WL [107]),
.WL108(WL [108]),
.WL109(WL [109]),
.WL110(WL [110]),
.WL111(WL [111]),
.WL112(WL [112]),
.WL113(WL [113]),
.WL114(WL [114]),
.WL115(WL [115]),
.WL116(WL [116]),
.WL117(WL [117]),
.WL118(WL [118]),
.WL119(WL [119]),
.WL120(WL [120]),
.WL121(WL [121]),
.WL122(WL [122]),
.WL123(WL [123]),
.WL124(WL [124]),
.WL125(WL [125]),
.WL126(WL [126]),
.WL127(WL [127]),
.WL128(WL [128]),
.WL129(WL [129]),
.WL130(WL [130]),
.WL131(WL [131]),
.WL132(WL [132]),
.WL133(WL [133]),
.WL134(WL [134]),
.WL135(WL [135]),
.WL136(WL [136]),
.WL137(WL [137]),
.WL138(WL [138]),
.WL139(WL [139]),
.WL140(WL [140]),
.WL141(WL [141]),
.WL142(WL [142]),
.WL143(WL [143]),
.WL144(WL [144]),
.WL145(WL [145]),
.WL146(WL [146]),
.WL147(WL [147]),
.WL148(WL [148]),
.WL149(WL [149]),
.WL150(WL [150]),
.WL151(WL [151]),
.WL152(WL [152]),
.WL153(WL [153]),
.WL154(WL [154]),
.WL155(WL [155]),
.WL156(WL [156]),
.WL157(WL [157]),
.WL158(WL [158]),
.WL159(WL [159]),
.WL160(WL [160]),
.WL161(WL [161]),
.WL162(WL [162]),
.WL163(WL [163]),
.WL164(WL [164]),
.WL165(WL [165]),
.WL166(WL [166]),
.WL167(WL [167]),
.WL168(WL [168]),
.WL169(WL [169]),
.WL170(WL [170]),
.WL171(WL [171]),
.WL172(WL [172]),
.WL173(WL [173]),
.WL174(WL [174]),
.WL175(WL [175]),
.WL176(WL [176]),
.WL177(WL [177]),
.WL178(WL [178]),
.WL179(WL [179]),
.WL180(WL [180]),
.WL181(WL [181]),
.WL182(WL [182]),
.WL183(WL [183]),
.WL184(WL [184]),
.WL185(WL [185]),
.WL186(WL [186]),
.WL187(WL [187]),
.WL188(WL [188]),
.WL189(WL [189]),
.WL190(WL [190]),
.WL191(WL [191]),
.WL192(WL [192]),
.WL193(WL [193]),
.WL194(WL [194]),
.WL195(WL [195]),
.WL196(WL [196]),
.WL197(WL [197]),
.WL198(WL [198]),
.WL199(WL [199]),
.WL200(WL [200]),
.WL201(WL [201]),
.WL202(WL [202]),
.WL203(WL [203]),
.WL204(WL [204]),
.WL205(WL [205]),
.WL206(WL [206]),
.WL207(WL [207]),
.WL208(WL [208]),
.WL209(WL [209]),
.WL210(WL [210]),
.WL211(WL [211]),
.WL212(WL [212]),
.WL213(WL [213]),
.WL214(WL [214]),
.WL215(WL [215]),
.WL216(WL [216]),
.WL217(WL [217]),
.WL218(WL [218]),
.WL219(WL [219]),
.WL220(WL [220]),
.WL221(WL [221]),
.WL222(WL [222]),
.WL223(WL [223]),
.WL224(WL [224]),
.WL225(WL [225]),
.WL226(WL [226]),
.WL227(WL [227]),
.WL228(WL [228]),
.WL229(WL [229]),
.WL230(WL [230]),
.WL231(WL [231]),
.WL232(WL [232]),
.WL233(WL [233]),
.WL234(WL [234]),
.WL235(WL [235]),
.WL236(WL [236]),
.WL237(WL [237]),
.WL238(WL [238]),
.WL239(WL [239]),
.WL240(WL [240]),
.WL241(WL [241]),
.WL242(WL [242]),
.WL243(WL [243]),
.WL244(WL [244]),
.WL245(WL [245]),
.WL246(WL [246]),
.WL247(WL [247]),
.WL248(WL [248]),
.WL249(WL [249]),
.WL250(WL [250]),
.WL251(WL [251]),
.WL252(WL [252]),
.WL253(WL [253]),
.WL254(WL [254]),
.WL255(WL [255]),
.WL256(WL [256]),
.WL257(WL [257]),
.WL258(WL [258]),
.WL259(WL [259]),
.WL260(WL [260]),
.WL261(WL [261]),
.WL262(WL [262]),
.WL263(WL [263]),
.WL264(WL [264]),
.WL265(WL [265]),
.WL266(WL [266]),
.WL267(WL [267]),
.WL268(WL [268]),
.WL269(WL [269]),
.WL270(WL [270]),
.WL271(WL [271]),
.WL272(WL [272]),
.WL273(WL [273]),
.WL274(WL [274]),
.WL275(WL [275]),
.WL276(WL [276]),
.WL277(WL [277]),
.WL278(WL [278]),
.WL279(WL [279]),
.WL280(WL [280]),
.WL281(WL [281]),
.WL282(WL [282]),
.WL283(WL [283]),
.WL284(WL [284]),
.WL285(WL [285]),
.WL286(WL [286]),
.WL287(WL [287]),
.WL288(WL [288]),
.WL289(WL [289]),
.WL290(WL [290]),
.WL291(WL [291]),
.WL292(WL [292]),
.WL293(WL [293]),
.WL294(WL [294]),
.WL295(WL [295]),
.WL296(WL [296]),
.WL297(WL [297]),
.WL298(WL [298]),
.WL299(WL [299]),
.WL300(WL [300]),
.WL301(WL [301]),
.WL302(WL [302]),
.WL303(WL [303]),
.WL304(WL [304]),
.WL305(WL [305]),
.WL306(WL [306]),
.WL307(WL [307]),
.WL308(WL [308]),
.WL309(WL [309]),
.WL310(WL [310]),
.WL311(WL [311]),
.WL312(WL [312]),
.WL313(WL [313]),
.WL314(WL [314]),
.WL315(WL [315]),
.WL316(WL [316]),
.WL317(WL [317]),
.WL318(WL [318]),
.WL319(WL [319]),
.WL320(WL [320]),
.WL321(WL [321]),
.WL322(WL [322]),
.WL323(WL [323]),
.WL324(WL [324]),
.WL325(WL [325]),
.WL326(WL [326]),
.WL327(WL [327]),
.WL328(WL [328]),
.WL329(WL [329]),
.WL330(WL [330]),
.WL331(WL [331]),
.WL332(WL [332]),
.WL333(WL [333]),
.WL334(WL [334]),
.WL335(WL [335]),
.WL336(WL [336]),
.WL337(WL [337]),
.WL338(WL [338]),
.WL339(WL [339]),
.WL340(WL [340]),
.WL341(WL [341]),
.WL342(WL [342]),
.WL343(WL [343]),
.WL344(WL [344]),
.WL345(WL [345]),
.WL346(WL [346]),
.WL347(WL [347]),
.WL348(WL [348]),
.WL349(WL [349]),
.WL350(WL [350]),
.WL351(WL [351]),
.WL352(WL [352]),
.WL353(WL [353]),
.WL354(WL [354]),
.WL355(WL [355]),
.WL356(WL [356]),
.WL357(WL [357]),
.WL358(WL [358]),
.WL359(WL [359]),
.WL360(WL [360]),
.WL361(WL [361]),
.WL362(WL [362]),
.WL363(WL [363]),
.WL364(WL [364]),
.WL365(WL [365]),
.WL366(WL [366]),
.WL367(WL [367]),
.WL368(WL [368]),
.WL369(WL [369]),
.WL370(WL [370]),
.WL371(WL [371]),
.WL372(WL [372]),
.WL373(WL [373]),
.WL374(WL [374]),
.WL375(WL [375]),
.WL376(WL [376]),
.WL377(WL [377]),
.WL378(WL [378]),
.WL379(WL [379]),
.WL380(WL [380]),
.WL381(WL [381]),
.WL382(WL [382]),
.WL383(WL [383]),
.WL384(WL [384]),
.WL385(WL [385]),
.WL386(WL [386]),
.WL387(WL [387]),
.WL388(WL [388]),
.WL389(WL [389]),
.WL390(WL [390]),
.WL391(WL [391]),
.WL392(WL [392]),
.WL393(WL [393]),
.WL394(WL [394]),
.WL395(WL [395]),
.WL396(WL [396]),
.WL397(WL [397]),
.WL398(WL [398]),
.WL399(WL [399]),
.WL400(WL [400]),
.WL401(WL [401]),
.WL402(WL [402]),
.WL403(WL [403]),
.WL404(WL [404]),
.WL405(WL [405]),
.WL406(WL [406]),
.WL407(WL [407]),
.WL408(WL [408]),
.WL409(WL [409]),
.WL410(WL [410]),
.WL411(WL [411]),
.WL412(WL [412]),
.WL413(WL [413]),
.WL414(WL [414]),
.WL415(WL [415]),
.WL416(WL [416]),
.WL417(WL [417]),
.WL418(WL [418]),
.WL419(WL [419]),
.WL420(WL [420]),
.WL421(WL [421]),
.WL422(WL [422]),
.WL423(WL [423]),
.WL424(WL [424]),
.WL425(WL [425]),
.WL426(WL [426]),
.WL427(WL [427]),
.WL428(WL [428]),
.WL429(WL [429]),
.WL430(WL [430]),
.WL431(WL [431]),
.WL432(WL [432]),
.WL433(WL [433]),
.WL434(WL [434]),
.WL435(WL [435]),
.WL436(WL [436]),
.WL437(WL [437]),
.WL438(WL [438]),
.WL439(WL [439]),
.WL440(WL [440]),
.WL441(WL [441]),
.WL442(WL [442]),
.WL443(WL [443]),
.WL444(WL [444]),
.WL445(WL [445]),
.WL446(WL [446]),
.WL447(WL [447]),
.WL448(WL [448]),
.WL449(WL [449]),
.WL450(WL [450]),
.WL451(WL [451]),
.WL452(WL [452]),
.WL453(WL [453]),
.WL454(WL [454]),
.WL455(WL [455]),
.WL456(WL [456]),
.WL457(WL [457]),
.WL458(WL [458]),
.WL459(WL [459]),
.WL460(WL [460]),
.WL461(WL [461]),
.WL462(WL [462]),
.WL463(WL [463]),
.WL464(WL [464]),
.WL465(WL [465]),
.WL466(WL [466]),
.WL467(WL [467]),
.WL468(WL [468]),
.WL469(WL [469]),
.WL470(WL [470]),
.WL471(WL [471]),
.WL472(WL [472]),
.WL473(WL [473]),
.WL474(WL [474]),
.WL475(WL [475]),
.WL476(WL [476]),
.WL477(WL [477]),
.WL478(WL [478]),
.WL479(WL [479]),
.WL480(WL [480]),
.WL481(WL [481]),
.WL482(WL [482]),
.WL483(WL [483]),
.WL484(WL [484]),
.WL485(WL [485]),
.WL486(WL [486]),
.WL487(WL [487]),
.WL488(WL [488]),
.WL489(WL [489]),
.WL490(WL [490]),
.WL491(WL [491]),
.WL492(WL [492]),
.WL493(WL [493]),
.WL494(WL [494]),
.WL495(WL [495]),
.WL496(WL [496]),
.WL497(WL [497]),
.WL498(WL [498]),
.WL499(WL [499]),
.WL500(WL [500]),
.WL501(WL [501]),
.WL502(WL [502]),
.WL503(WL [503]),
.WL504(WL [504]),
.WL505(WL [505]),
.WL506(WL [506]),
.WL507(WL [507]),
.WL508(WL [508]),
.WL509(WL [509]),
.WL510(WL [510]),
.WL511(WL [511]),
.WL512(WL [512]),
.WL513(WL [513]),
.WL514(WL [514]),
.WL515(WL [515]),
.WL516(WL [516]),
.WL517(WL [517]),
.WL518(WL [518]),
.WL519(WL [519]),
.WL520(WL [520]),
.WL521(WL [521]),
.WL522(WL [522]),
.WL523(WL [523]),
.WL524(WL [524]),
.WL525(WL [525]),
.WL526(WL [526]),
.WL527(WL [527]),
.WL528(WL [528]),
.WL529(WL [529]),
.WL530(WL [530]),
.WL531(WL [531]),
.WL532(WL [532]),
.WL533(WL [533]),
.WL534(WL [534]),
.WL535(WL [535]),
.WL536(WL [536]),
.WL537(WL [537]),
.WL538(WL [538]),
.WL539(WL [539]),
.WL540(WL [540]),
.WL541(WL [541]),
.WL542(WL [542]),
.WL543(WL [543]),
.WL544(WL [544]),
.WL545(WL [545]),
.WL546(WL [546]),
.WL547(WL [547]),
.WL548(WL [548]),
.WL549(WL [549]),
.WL550(WL [550]),
.WL551(WL [551]),
.WL552(WL [552]),
.WL553(WL [553]),
.WL554(WL [554]),
.WL555(WL [555]),
.WL556(WL [556]),
.WL557(WL [557]),
.WL558(WL [558]),
.WL559(WL [559]),
.WL560(WL [560]),
.WL561(WL [561]),
.WL562(WL [562]),
.WL563(WL [563]),
.WL564(WL [564]),
.WL565(WL [565]),
.WL566(WL [566]),
.WL567(WL [567]),
.WL568(WL [568]),
.WL569(WL [569]),
.WL570(WL [570]),
.WL571(WL [571]),
.WL572(WL [572]),
.WL573(WL [573]),
.WL574(WL [574]),
.WL575(WL [575]),
.WL576(WL [576]),
.WL577(WL [577]),
.WL578(WL [578]),
.WL579(WL [579]),
.WL580(WL [580]),
.WL581(WL [581]),
.WL582(WL [582]),
.WL583(WL [583]),
.WL584(WL [584]),
.WL585(WL [585]),
.WL586(WL [586]),
.WL587(WL [587]),
.WL588(WL [588]),
.WL589(WL [589]),
.WL590(WL [590]),
.WL591(WL [591]),
.WL592(WL [592]),
.WL593(WL [593]),
.WL594(WL [594]),
.WL595(WL [595]),
.WL596(WL [596]),
.WL597(WL [597]),
.WL598(WL [598]),
.WL599(WL [599]),
.WL600(WL [600]),
.WL601(WL [601]),
.WL602(WL [602]),
.WL603(WL [603]),
.WL604(WL [604]),
.WL605(WL [605]),
.WL606(WL [606]),
.WL607(WL [607]),
.WL608(WL [608]),
.WL609(WL [609]),
.WL610(WL [610]),
.WL611(WL [611]),
.WL612(WL [612]),
.WL613(WL [613]),
.WL614(WL [614]),
.WL615(WL [615]),
.WL616(WL [616]),
.WL617(WL [617]),
.WL618(WL [618]),
.WL619(WL [619]),
.WL620(WL [620]),
.WL621(WL [621]),
.WL622(WL [622]),
.WL623(WL [623]),
.WL624(WL [624]),
.WL625(WL [625]),
.WL626(WL [626]),
.WL627(WL [627]),
.WL628(WL [628]),
.WL629(WL [629]),
.WL630(WL [630]),
.WL631(WL [631]),
.WL632(WL [632]),
.WL633(WL [633]),
.WL634(WL [634]),
.WL635(WL [635]),
.WL636(WL [636]),
.WL637(WL [637]),
.WL638(WL [638]),
.WL639(WL [639]),
.WL640(WL [640]),
.WL641(WL [641]),
.WL642(WL [642]),
.WL643(WL [643]),
.WL644(WL [644]),
.WL645(WL [645]),
.WL646(WL [646]),
.WL647(WL [647]),
.WL648(WL [648]),
.WL649(WL [649]),
.WL650(WL [650]),
.WL651(WL [651]),
.WL652(WL [652]),
.WL653(WL [653]),
.WL654(WL [654]),
.WL655(WL [655]),
.WL656(WL [656]),
.WL657(WL [657]),
.WL658(WL [658]),
.WL659(WL [659]),
.WL660(WL [660]),
.WL661(WL [661]),
.WL662(WL [662]),
.WL663(WL [663]),
.WL664(WL [664]),
.WL665(WL [665]),
.WL666(WL [666]),
.WL667(WL [667]),
.WL668(WL [668]),
.WL669(WL [669]),
.WL670(WL [670]),
.WL671(WL [671]),
.WL672(WL [672]),
.WL673(WL [673]),
.WL674(WL [674]),
.WL675(WL [675]),
.WL676(WL [676]),
.WL677(WL [677]),
.WL678(WL [678]),
.WL679(WL [679]),
.WL680(WL [680]),
.WL681(WL [681]),
.WL682(WL [682]),
.WL683(WL [683]),
.WL684(WL [684]),
.WL685(WL [685]),
.WL686(WL [686]),
.WL687(WL [687]),
.WL688(WL [688]),
.WL689(WL [689]),
.WL690(WL [690]),
.WL691(WL [691]),
.WL692(WL [692]),
.WL693(WL [693]),
.WL694(WL [694]),
.WL695(WL [695]),
.WL696(WL [696]),
.WL697(WL [697]),
.WL698(WL [698]),
.WL699(WL [699]),
.WL700(WL [700]),
.WL701(WL [701]),
.WL702(WL [702]),
.WL703(WL [703]),
.WL704(WL [704]),
.WL705(WL [705]),
.WL706(WL [706]),
.WL707(WL [707]),
.WL708(WL [708]),
.WL709(WL [709]),
.WL710(WL [710]),
.WL711(WL [711]),
.WL712(WL [712]),
.WL713(WL [713]),
.WL714(WL [714]),
.WL715(WL [715]),
.WL716(WL [716]),
.WL717(WL [717]),
.WL718(WL [718]),
.WL719(WL [719]),
.WL720(WL [720]),
.WL721(WL [721]),
.WL722(WL [722]),
.WL723(WL [723]),
.WL724(WL [724]),
.WL725(WL [725]),
.WL726(WL [726]),
.WL727(WL [727]),
.WL728(WL [728]),
.WL729(WL [729]),
.WL730(WL [730]),
.WL731(WL [731]),
.WL732(WL [732]),
.WL733(WL [733]),
.WL734(WL [734]),
.WL735(WL [735]),
.WL736(WL [736]),
.WL737(WL [737]),
.WL738(WL [738]),
.WL739(WL [739]),
.WL740(WL [740]),
.WL741(WL [741]),
.WL742(WL [742]),
.WL743(WL [743]),
.WL744(WL [744]),
.WL745(WL [745]),
.WL746(WL [746]),
.WL747(WL [747]),
.WL748(WL [748]),
.WL749(WL [749]),
.WL750(WL [750]),
.WL751(WL [751]),
.WL752(WL [752]),
.WL753(WL [753]),
.WL754(WL [754]),
.WL755(WL [755]),
.WL756(WL [756]),
.WL757(WL [757]),
.WL758(WL [758]),
.WL759(WL [759]),
.WL760(WL [760]),
.WL761(WL [761]),
.WL762(WL [762]),
.WL763(WL [763]),
.WL764(WL [764]),
.WL765(WL [765]),
.WL766(WL [766]),
.WL767(WL [767]),
.WL768(WL [768]),
.WL769(WL [769]),
.WL770(WL [770]),
.WL771(WL [771]),
.WL772(WL [772]),
.WL773(WL [773]),
.WL774(WL [774]),
.WL775(WL [775]),
.WL776(WL [776]),
.WL777(WL [777]),
.WL778(WL [778]),
.WL779(WL [779]),
.WL780(WL [780]),
.WL781(WL [781]),
.WL782(WL [782]),
.WL783(WL [783]),
.WL784(WL [784]),
.WL785(WL [785]),
.WL786(WL [786]),
.WL787(WL [787]),
.WL788(WL [788]),
.WL789(WL [789]),
.WL790(WL [790]),
.WL791(WL [791]),
.WL792(WL [792]),
.WL793(WL [793]),
.WL794(WL [794]),
.WL795(WL [795]),
.WL796(WL [796]),
.WL797(WL [797]),
.WL798(WL [798]),
.WL799(WL [799]),
.WL800(WL [800]),
.WL801(WL [801]),
.WL802(WL [802]),
.WL803(WL [803]),
.WL804(WL [804]),
.WL805(WL [805]),
.WL806(WL [806]),
.WL807(WL [807]),
.WL808(WL [808]),
.WL809(WL [809]),
.WL810(WL [810]),
.WL811(WL [811]),
.WL812(WL [812]),
.WL813(WL [813]),
.WL814(WL [814]),
.WL815(WL [815]),
.WL816(WL [816]),
.WL817(WL [817]),
.WL818(WL [818]),
.WL819(WL [819]),
.WL820(WL [820]),
.WL821(WL [821]),
.WL822(WL [822]),
.WL823(WL [823]),
.WL824(WL [824]),
.WL825(WL [825]),
.WL826(WL [826]),
.WL827(WL [827]),
.WL828(WL [828]),
.WL829(WL [829]),
.WL830(WL [830]),
.WL831(WL [831]),
.WL832(WL [832]),
.WL833(WL [833]),
.WL834(WL [834]),
.WL835(WL [835]),
.WL836(WL [836]),
.WL837(WL [837]),
.WL838(WL [838]),
.WL839(WL [839]),
.WL840(WL [840]),
.WL841(WL [841]),
.WL842(WL [842]),
.WL843(WL [843]),
.WL844(WL [844]),
.WL845(WL [845]),
.WL846(WL [846]),
.WL847(WL [847]),
.WL848(WL [848]),
.WL849(WL [849]),
.WL850(WL [850]),
.WL851(WL [851]),
.WL852(WL [852]),
.WL853(WL [853]),
.WL854(WL [854]),
.WL855(WL [855]),
.WL856(WL [856]),
.WL857(WL [857]),
.WL858(WL [858]),
.WL859(WL [859]),
.WL860(WL [860]),
.WL861(WL [861]),
.WL862(WL [862]),
.WL863(WL [863]),
.WL864(WL [864]),
.WL865(WL [865]),
.WL866(WL [866]),
.WL867(WL [867]),
.WL868(WL [868]),
.WL869(WL [869]),
.WL870(WL [870]),
.WL871(WL [871]),
.WL872(WL [872]),
.WL873(WL [873]),
.WL874(WL [874]),
.WL875(WL [875]),
.WL876(WL [876]),
.WL877(WL [877]),
.WL878(WL [878]),
.WL879(WL [879]),
.WL880(WL [880]),
.WL881(WL [881]),
.WL882(WL [882]),
.WL883(WL [883]),
.WL884(WL [884]),
.WL885(WL [885]),
.WL886(WL [886]),
.WL887(WL [887]),
.WL888(WL [888]),
.WL889(WL [889]),
.WL890(WL [890]),
.WL891(WL [891]),
.WL892(WL [892]),
.WL893(WL [893]),
.WL894(WL [894]),
.WL895(WL [895]),
.WL896(WL [896]),
.WL897(WL [897]),
.WL898(WL [898]),
.WL899(WL [899]),
.WL900(WL [900]),
.WL901(WL [901]),
.WL902(WL [902]),
.WL903(WL [903]),
.WL904(WL [904]),
.WL905(WL [905]),
.WL906(WL [906]),
.WL907(WL [907]),
.WL908(WL [908]),
.WL909(WL [909]),
.WL910(WL [910]),
.WL911(WL [911]),
.WL912(WL [912]),
.WL913(WL [913]),
.WL914(WL [914]),
.WL915(WL [915]),
.WL916(WL [916]),
.WL917(WL [917]),
.WL918(WL [918]),
.WL919(WL [919]),
.WL920(WL [920]),
.WL921(WL [921]),
.WL922(WL [922]),
.WL923(WL [923]),
.WL924(WL [924]),
.WL925(WL [925]),
.WL926(WL [926]),
.WL927(WL [927]),
.WL928(WL [928]),
.WL929(WL [929]),
.WL930(WL [930]),
.WL931(WL [931]),
.WL932(WL [932]),
.WL933(WL [933]),
.WL934(WL [934]),
.WL935(WL [935]),
.WL936(WL [936]),
.WL937(WL [937]),
.WL938(WL [938]),
.WL939(WL [939]),
.WL940(WL [940]),
.WL941(WL [941]),
.WL942(WL [942]),
.WL943(WL [943]),
.WL944(WL [944]),
.WL945(WL [945]),
.WL946(WL [946]),
.WL947(WL [947]),
.WL948(WL [948]),
.WL949(WL [949]),
.WL950(WL [950]),
.WL951(WL [951]),
.WL952(WL [952]),
.WL953(WL [953]),
.WL954(WL [954]),
.WL955(WL [955]),
.WL956(WL [956]),
.WL957(WL [957]),
.WL958(WL [958]),
.WL959(WL [959]),
.WL960(WL [960]),
.WL961(WL [961]),
.WL962(WL [962]),
.WL963(WL [963]),
.WL964(WL [964]),
.WL965(WL [965]),
.WL966(WL [966]),
.WL967(WL [967]),
.WL968(WL [968]),
.WL969(WL [969]),
.WL970(WL [970]),
.WL971(WL [971]),
.WL972(WL [972]),
.WL973(WL [973]),
.WL974(WL [974]),
.WL975(WL [975]),
.WL976(WL [976]),
.WL977(WL [977]),
.WL978(WL [978]),
.WL979(WL [979]),
.WL980(WL [980]),
.WL981(WL [981]),
.WL982(WL [982]),
.WL983(WL [983]),
.WL984(WL [984]),
.WL985(WL [985]),
.WL986(WL [986]),
.WL987(WL [987]),
.WL988(WL [988]),
.WL989(WL [989]),
.WL990(WL [990]),
.WL991(WL [991]),
.WL992(WL [992]),
.WL993(WL [993]),
.WL994(WL [994]),
.WL995(WL [995]),
.WL996(WL [996]),
.WL997(WL [997]),
.WL998(WL [998]),
.WL999(WL [999]),
.WL1000(WL [1000]),
.WL1001(WL [1001]),
.WL1002(WL [1002]),
.WL1003(WL [1003]),
.WL1004(WL [1004]),
.WL1005(WL [1005]),
.WL1006(WL [1006]),
.WL1007(WL [1007]),
.WL1008(WL [1008]),
.WL1009(WL [1009]),
.WL1010(WL [1010]),
.WL1011(WL [1011]),
.WL1012(WL [1012]),
.WL1013(WL [1013]),
.WL1014(WL [1014]),
.WL1015(WL [1015]),
.WL1016(WL [1016]),
.WL1017(WL [1017]),
.WL1018(WL [1018]),
.WL1019(WL [1019]),
.WL1020(WL [1020]),
.WL1021(WL [1021]),
.WL1022(WL [1022]),
.WL1023(WL [1023])

);



endmodule








