VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO IMPACTSram
  CLASS BLOCK ;
  FOREIGN IMPACTSram ;
  ORIGIN 3.500 45.700 ;
  SIZE 236.200 BY 68.000 ;
  PIN BL0
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met2 ;
        RECT 1.500 22.000 1.800 22.300 ;
    END
  END BL0
  PIN BLb0
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met2 ;
        RECT 6.600 22.000 6.900 22.300 ;
    END
  END BLb0
  PIN BLb1
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met2 ;
        RECT 13.350 22.000 13.650 22.300 ;
    END
  END BLb1
  PIN BL31
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met2 ;
        RECT 210.750 22.000 211.050 22.300 ;
    END
  END BL31
  PIN BL30
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met2 ;
        RECT 204.000 22.000 204.300 22.300 ;
    END
  END BL30
  PIN BL29
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met2 ;
        RECT 197.250 22.000 197.550 22.300 ;
    END
  END BL29
  PIN BL28
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met2 ;
        RECT 190.500 22.000 190.800 22.300 ;
    END
  END BL28
  PIN BL27
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met2 ;
        RECT 183.750 22.000 184.050 22.300 ;
    END
  END BL27
  PIN BL26
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met2 ;
        RECT 177.000 22.000 177.300 22.300 ;
    END
  END BL26
  PIN BL25
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met2 ;
        RECT 170.250 22.000 170.550 22.300 ;
    END
  END BL25
  PIN BL24
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met2 ;
        RECT 163.500 22.000 163.800 22.300 ;
    END
  END BL24
  PIN BL23
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met2 ;
        RECT 156.800 22.000 157.100 22.300 ;
    END
  END BL23
  PIN BL22
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met2 ;
        RECT 150.000 22.000 150.300 22.300 ;
    END
  END BL22
  PIN BL21
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met2 ;
        RECT 143.250 22.000 143.550 22.300 ;
    END
  END BL21
  PIN BL20
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met2 ;
        RECT 136.500 22.000 136.800 22.300 ;
    END
  END BL20
  PIN BL19
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met2 ;
        RECT 129.750 22.000 130.050 22.300 ;
    END
  END BL19
  PIN BL18
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met2 ;
        RECT 123.000 22.000 123.300 22.300 ;
    END
  END BL18
  PIN BL17
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met2 ;
        RECT 116.250 22.000 116.550 22.300 ;
    END
  END BL17
  PIN BL16
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met2 ;
        RECT 109.500 22.000 109.800 22.300 ;
    END
  END BL16
  PIN BL15
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met2 ;
        RECT 102.750 22.000 103.050 22.300 ;
    END
  END BL15
  PIN BL14
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met2 ;
        RECT 96.000 22.000 96.300 22.300 ;
    END
  END BL14
  PIN BL13
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met2 ;
        RECT 89.250 22.000 89.550 22.300 ;
    END
  END BL13
  PIN BL12
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met2 ;
        RECT 82.500 22.000 82.800 22.300 ;
    END
  END BL12
  PIN BL11
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met2 ;
        RECT 75.750 22.000 76.050 22.300 ;
    END
  END BL11
  PIN BL10
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met2 ;
        RECT 69.000 22.000 69.300 22.300 ;
    END
  END BL10
  PIN BL9
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met2 ;
        RECT 62.250 22.000 62.550 22.300 ;
    END
  END BL9
  PIN BL8
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met2 ;
        RECT 55.500 22.000 55.800 22.300 ;
    END
  END BL8
  PIN BL7
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met2 ;
        RECT 48.750 22.000 49.050 22.300 ;
    END
  END BL7
  PIN BL6
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met2 ;
        RECT 42.000 22.000 42.300 22.300 ;
    END
  END BL6
  PIN BL5
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met2 ;
        RECT 35.250 22.000 35.550 22.300 ;
    END
  END BL5
  PIN BL4
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met2 ;
        RECT 28.500 22.000 28.800 22.300 ;
    END
  END BL4
  PIN BL3
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met2 ;
        RECT 21.750 22.000 22.050 22.300 ;
    END
  END BL3
  PIN BL2
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met2 ;
        RECT 15.000 22.000 15.300 22.300 ;
    END
  END BL2
  PIN BL1
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met2 ;
        RECT 8.200 22.000 8.500 22.300 ;
    END
  END BL1
  PIN BLb2
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met2 ;
        RECT 20.100 22.000 20.400 22.300 ;
    END
  END BLb2
  PIN BLb3
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met2 ;
        RECT 26.850 22.000 27.150 22.300 ;
    END
  END BLb3
  PIN BLb4
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met2 ;
        RECT 33.600 22.000 33.900 22.300 ;
    END
  END BLb4
  PIN BLb5
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met2 ;
        RECT 40.350 22.000 40.650 22.300 ;
    END
  END BLb5
  PIN BLb6
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met2 ;
        RECT 47.100 22.000 47.400 22.300 ;
    END
  END BLb6
  PIN BLb7
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met2 ;
        RECT 53.850 22.000 54.150 22.300 ;
    END
  END BLb7
  PIN BLb8
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met2 ;
        RECT 60.600 22.000 60.900 22.300 ;
    END
  END BLb8
  PIN BLb9
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met2 ;
        RECT 67.350 22.000 67.650 22.300 ;
    END
  END BLb9
  PIN BLb10
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met2 ;
        RECT 74.100 22.000 74.400 22.300 ;
    END
  END BLb10
  PIN BLb11
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met2 ;
        RECT 80.850 22.000 81.150 22.300 ;
    END
  END BLb11
  PIN BLb12
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met2 ;
        RECT 87.550 22.000 87.850 22.300 ;
    END
  END BLb12
  PIN BLb13
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met2 ;
        RECT 94.300 22.000 94.600 22.300 ;
    END
  END BLb13
  PIN BLb14
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met2 ;
        RECT 101.050 22.000 101.350 22.300 ;
    END
  END BLb14
  PIN BLb15
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met2 ;
        RECT 107.800 22.000 108.100 22.300 ;
    END
  END BLb15
  PIN BLb16
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met2 ;
        RECT 114.600 22.000 114.900 22.300 ;
    END
  END BLb16
  PIN BLb17
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met2 ;
        RECT 121.300 22.000 121.600 22.300 ;
    END
  END BLb17
  PIN BLb18
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met2 ;
        RECT 128.050 22.000 128.350 22.300 ;
    END
  END BLb18
  PIN BLb19
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met2 ;
        RECT 134.850 22.000 135.150 22.300 ;
    END
  END BLb19
  PIN BLb20
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met2 ;
        RECT 141.600 22.000 141.900 22.300 ;
    END
  END BLb20
  PIN BLb21
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met2 ;
        RECT 148.350 22.000 148.650 22.300 ;
    END
  END BLb21
  PIN BLb22
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met2 ;
        RECT 155.150 22.000 155.450 22.300 ;
    END
  END BLb22
  PIN BLb23
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met2 ;
        RECT 161.800 22.000 162.100 22.300 ;
    END
  END BLb23
  PIN BLb24
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met2 ;
        RECT 168.600 22.000 168.900 22.300 ;
    END
  END BLb24
  PIN BLb25
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met2 ;
        RECT 175.350 22.000 175.650 22.300 ;
    END
  END BLb25
  PIN BLb26
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met2 ;
        RECT 182.100 22.000 182.400 22.300 ;
    END
  END BLb26
  PIN BLb27
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met2 ;
        RECT 188.800 22.000 189.100 22.300 ;
    END
  END BLb27
  PIN BLb28
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met2 ;
        RECT 195.600 22.000 195.900 22.300 ;
    END
  END BLb28
  PIN BLb29
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met2 ;
        RECT 202.350 22.000 202.650 22.300 ;
    END
  END BLb29
  PIN BLb30
    ANTENNADIFFAREA 6.569000 ;
    PORT
      LAYER met2 ;
        RECT 209.100 22.000 209.400 22.300 ;
    END
  END BLb30
  PIN BLb31
    ANTENNADIFFAREA 6.184000 ;
    PORT
      LAYER met2 ;
        RECT 215.850 22.000 216.150 22.300 ;
    END
  END BLb31
  PIN WL0
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER met3 ;
        RECT -3.500 15.700 -2.900 16.300 ;
    END
  END WL0
  PIN WL1
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER met3 ;
        RECT -3.500 13.850 -2.900 14.450 ;
    END
  END WL1
  PIN WL2
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER met3 ;
        RECT -3.500 12.100 -2.900 12.700 ;
    END
  END WL2
  PIN WL3
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER met3 ;
        RECT -3.500 10.250 -2.900 10.850 ;
    END
  END WL3
  PIN WL4
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER met3 ;
        RECT -3.500 8.450 -2.900 9.050 ;
    END
  END WL4
  PIN WL5
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER met3 ;
        RECT -3.500 6.600 -2.900 7.200 ;
    END
  END WL5
  PIN WL6
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER met3 ;
        RECT -3.500 4.850 -2.900 5.450 ;
    END
  END WL6
  PIN WL7
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER met3 ;
        RECT -3.500 3.000 -2.900 3.600 ;
    END
  END WL7
  PIN WL8
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER met3 ;
        RECT -3.500 1.250 -2.900 1.850 ;
    END
  END WL8
  PIN WL9
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER met3 ;
        RECT -3.500 -0.600 -2.900 0.000 ;
    END
  END WL9
  PIN WL10
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER met3 ;
        RECT -3.500 -2.350 -2.900 -1.750 ;
    END
  END WL10
  PIN WL11
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER met3 ;
        RECT -3.500 -4.200 -2.900 -3.600 ;
    END
  END WL11
  PIN WL12
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER met3 ;
        RECT -3.500 -6.000 -2.900 -5.400 ;
    END
  END WL12
  PIN WL13
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER met3 ;
        RECT -3.500 -7.850 -2.900 -7.250 ;
    END
  END WL13
  PIN WL14
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER met3 ;
        RECT -3.500 -9.600 -2.900 -9.000 ;
    END
  END WL14
  PIN WL15
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER met3 ;
        RECT -3.500 -11.450 -2.900 -10.850 ;
    END
  END WL15
  PIN WL16
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER met3 ;
        RECT -3.500 -13.200 -2.900 -12.600 ;
    END
  END WL16
  PIN WL17
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER met3 ;
        RECT -3.500 -15.050 -2.900 -14.450 ;
    END
  END WL17
  PIN WL18
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER met3 ;
        RECT -3.500 -16.800 -2.900 -16.200 ;
    END
  END WL18
  PIN WL19
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER met3 ;
        RECT -3.500 -18.650 -2.900 -18.050 ;
    END
  END WL19
  PIN WL20
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER met3 ;
        RECT -3.500 -20.450 -2.900 -19.850 ;
    END
  END WL20
  PIN WL21
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER met3 ;
        RECT -3.500 -22.300 -2.900 -21.700 ;
    END
  END WL21
  PIN WL22
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER met3 ;
        RECT -3.500 -24.050 -2.900 -23.450 ;
    END
  END WL22
  PIN WL23
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER met3 ;
        RECT -3.500 -25.900 -2.900 -25.300 ;
    END
  END WL23
  PIN WL24
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER met3 ;
        RECT -3.500 -27.600 -2.900 -27.000 ;
    END
  END WL24
  PIN WL25
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER met3 ;
        RECT -3.500 -29.450 -2.900 -28.850 ;
    END
  END WL25
  PIN WL26
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER met3 ;
        RECT -3.500 -31.200 -2.900 -30.600 ;
    END
  END WL26
  PIN WL27
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER met3 ;
        RECT -3.500 -33.050 -2.900 -32.450 ;
    END
  END WL27
  PIN WL28
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER met3 ;
        RECT -3.500 -34.850 -2.900 -34.250 ;
    END
  END WL28
  PIN WL29
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER met3 ;
        RECT -3.500 -36.700 -2.900 -36.100 ;
    END
  END WL29
  PIN WL30
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER met3 ;
        RECT -3.500 -38.450 -2.900 -37.850 ;
    END
  END WL30
  PIN WL31
    ANTENNAGATEAREA 4.032000 ;
    PORT
      LAYER met3 ;
        RECT -3.500 -40.300 -2.900 -39.700 ;
    END
  END WL31
  PIN vccd1
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT -3.500 21.100 232.700 21.700 ;
    END
  END vccd1
  PIN vssd1
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT -3.500 19.400 232.700 19.900 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT -1.100 -41.100 218.900 17.120 ;
      LAYER met1 ;
        RECT -1.100 -43.350 218.900 22.300 ;
      LAYER met2 ;
        RECT -2.900 21.720 1.220 22.300 ;
        RECT 2.080 21.720 6.320 22.300 ;
        RECT 7.180 21.720 7.920 22.300 ;
        RECT 8.780 21.720 13.070 22.300 ;
        RECT 13.930 21.720 14.720 22.300 ;
        RECT 15.580 21.720 19.820 22.300 ;
        RECT 20.680 21.720 21.470 22.300 ;
        RECT 22.330 21.720 26.570 22.300 ;
        RECT 27.430 21.720 28.220 22.300 ;
        RECT 29.080 21.720 33.320 22.300 ;
        RECT 34.180 21.720 34.970 22.300 ;
        RECT 35.830 21.720 40.070 22.300 ;
        RECT 40.930 21.720 41.720 22.300 ;
        RECT 42.580 21.720 46.820 22.300 ;
        RECT 47.680 21.720 48.470 22.300 ;
        RECT 49.330 21.720 53.570 22.300 ;
        RECT 54.430 21.720 55.220 22.300 ;
        RECT 56.080 21.720 60.320 22.300 ;
        RECT 61.180 21.720 61.970 22.300 ;
        RECT 62.830 21.720 67.070 22.300 ;
        RECT 67.930 21.720 68.720 22.300 ;
        RECT 69.580 21.720 73.820 22.300 ;
        RECT 74.680 21.720 75.470 22.300 ;
        RECT 76.330 21.720 80.570 22.300 ;
        RECT 81.430 21.720 82.220 22.300 ;
        RECT 83.080 21.720 87.270 22.300 ;
        RECT 88.130 21.720 88.970 22.300 ;
        RECT 89.830 21.720 94.020 22.300 ;
        RECT 94.880 21.720 95.720 22.300 ;
        RECT 96.580 21.720 100.770 22.300 ;
        RECT 101.630 21.720 102.470 22.300 ;
        RECT 103.330 21.720 107.520 22.300 ;
        RECT 108.380 21.720 109.220 22.300 ;
        RECT 110.080 21.720 114.320 22.300 ;
        RECT 115.180 21.720 115.970 22.300 ;
        RECT 116.830 21.720 121.020 22.300 ;
        RECT 121.880 21.720 122.720 22.300 ;
        RECT 123.580 21.720 127.770 22.300 ;
        RECT 128.630 21.720 129.470 22.300 ;
        RECT 130.330 21.720 134.570 22.300 ;
        RECT 135.430 21.720 136.220 22.300 ;
        RECT 137.080 21.720 141.320 22.300 ;
        RECT 142.180 21.720 142.970 22.300 ;
        RECT 143.830 21.720 148.070 22.300 ;
        RECT 148.930 21.720 149.720 22.300 ;
        RECT 150.580 21.720 154.870 22.300 ;
        RECT 155.730 21.720 156.520 22.300 ;
        RECT 157.380 21.720 161.520 22.300 ;
        RECT 162.380 21.720 163.220 22.300 ;
        RECT 164.080 21.720 168.320 22.300 ;
        RECT 169.180 21.720 169.970 22.300 ;
        RECT 170.830 21.720 175.070 22.300 ;
        RECT 175.930 21.720 176.720 22.300 ;
        RECT 177.580 21.720 181.820 22.300 ;
        RECT 182.680 21.720 183.470 22.300 ;
        RECT 184.330 21.720 188.520 22.300 ;
        RECT 189.380 21.720 190.220 22.300 ;
        RECT 191.080 21.720 195.320 22.300 ;
        RECT 196.180 21.720 196.970 22.300 ;
        RECT 197.830 21.720 202.070 22.300 ;
        RECT 202.930 21.720 203.720 22.300 ;
        RECT 204.580 21.720 208.820 22.300 ;
        RECT 209.680 21.720 210.470 22.300 ;
        RECT 211.330 21.720 215.570 22.300 ;
        RECT 216.430 21.720 220.700 22.300 ;
        RECT -2.900 -45.700 220.700 21.720 ;
      LAYER met3 ;
        RECT -3.500 16.300 -2.900 16.600 ;
        RECT -3.500 15.400 -2.900 15.700 ;
        RECT -2.500 15.300 220.700 16.600 ;
        RECT -3.500 14.850 220.700 15.300 ;
        RECT -3.500 14.450 -2.900 14.750 ;
        RECT -3.500 13.550 -2.900 13.850 ;
        RECT -2.500 13.450 220.700 14.850 ;
        RECT -3.500 13.100 220.700 13.450 ;
        RECT -3.500 12.700 -2.900 13.000 ;
        RECT -3.500 11.800 -2.900 12.100 ;
        RECT -2.500 11.700 220.700 13.100 ;
        RECT -3.500 11.250 220.700 11.700 ;
        RECT -3.500 10.850 -2.900 11.150 ;
        RECT -3.500 9.950 -2.900 10.250 ;
        RECT -2.500 9.850 220.700 11.250 ;
        RECT -3.500 9.450 220.700 9.850 ;
        RECT -3.500 9.050 -2.900 9.350 ;
        RECT -3.500 8.150 -2.900 8.450 ;
        RECT -2.500 8.050 220.700 9.450 ;
        RECT -3.500 7.600 220.700 8.050 ;
        RECT -3.500 7.200 -2.900 7.500 ;
        RECT -3.500 6.300 -2.900 6.600 ;
        RECT -2.500 6.200 220.700 7.600 ;
        RECT -3.500 5.850 220.700 6.200 ;
        RECT -3.500 5.450 -2.900 5.750 ;
        RECT -3.500 4.550 -2.900 4.850 ;
        RECT -2.500 4.450 220.700 5.850 ;
        RECT -3.500 4.000 220.700 4.450 ;
        RECT -3.500 3.600 -2.900 3.900 ;
        RECT -3.500 2.700 -2.900 3.000 ;
        RECT -2.500 2.600 220.700 4.000 ;
        RECT -3.500 2.250 220.700 2.600 ;
        RECT -3.500 1.850 -2.900 2.150 ;
        RECT -3.500 0.950 -2.900 1.250 ;
        RECT -2.500 0.850 220.700 2.250 ;
        RECT -3.500 0.400 220.700 0.850 ;
        RECT -3.500 0.000 -2.900 0.300 ;
        RECT -3.500 -0.900 -2.900 -0.600 ;
        RECT -2.500 -1.000 220.700 0.400 ;
        RECT -3.500 -1.350 220.700 -1.000 ;
        RECT -3.500 -1.750 -2.900 -1.400 ;
        RECT -3.500 -2.600 -2.900 -2.350 ;
        RECT -2.500 -2.750 220.700 -1.350 ;
        RECT -3.500 -3.200 220.700 -2.750 ;
        RECT -3.500 -3.600 -2.900 -3.300 ;
        RECT -3.500 -4.500 -2.900 -4.200 ;
        RECT -2.500 -4.600 220.700 -3.200 ;
        RECT -3.500 -5.000 220.700 -4.600 ;
        RECT -3.500 -5.400 -2.900 -5.100 ;
        RECT -3.500 -6.300 -2.900 -6.000 ;
        RECT -2.500 -6.400 220.700 -5.000 ;
        RECT -3.500 -6.850 220.700 -6.400 ;
        RECT -3.500 -7.250 -2.900 -6.900 ;
        RECT -3.500 -8.100 -2.900 -7.850 ;
        RECT -2.500 -8.250 220.700 -6.850 ;
        RECT -3.500 -8.600 220.700 -8.250 ;
        RECT -3.500 -9.000 -2.900 -8.700 ;
        RECT -3.500 -9.900 -2.900 -9.600 ;
        RECT -2.500 -10.000 220.700 -8.600 ;
        RECT -3.500 -10.450 220.700 -10.000 ;
        RECT -3.500 -10.850 -2.900 -10.500 ;
        RECT -3.500 -11.700 -2.900 -11.450 ;
        RECT -2.500 -11.850 220.700 -10.450 ;
        RECT -3.500 -12.200 220.700 -11.850 ;
        RECT -3.500 -12.600 -2.900 -12.300 ;
        RECT -3.500 -13.500 -2.900 -13.200 ;
        RECT -2.500 -13.600 220.700 -12.200 ;
        RECT -3.500 -14.050 220.700 -13.600 ;
        RECT -3.500 -14.450 -2.900 -14.100 ;
        RECT -3.500 -15.300 -2.900 -15.050 ;
        RECT -2.500 -15.450 220.700 -14.050 ;
        RECT -3.500 -15.800 220.700 -15.450 ;
        RECT -3.500 -16.200 -2.900 -15.900 ;
        RECT -3.500 -17.100 -2.900 -16.800 ;
        RECT -2.500 -17.200 220.700 -15.800 ;
        RECT -3.500 -17.650 220.700 -17.200 ;
        RECT -3.500 -18.050 -2.900 -17.700 ;
        RECT -3.500 -18.900 -2.900 -18.650 ;
        RECT -2.500 -19.050 220.700 -17.650 ;
        RECT -3.500 -19.450 220.700 -19.050 ;
        RECT -3.500 -19.850 -2.900 -19.500 ;
        RECT -3.500 -20.700 -2.900 -20.450 ;
        RECT -2.500 -20.850 220.700 -19.450 ;
        RECT -3.500 -21.300 220.700 -20.850 ;
        RECT -3.500 -21.700 -2.900 -21.400 ;
        RECT -3.500 -22.600 -2.900 -22.300 ;
        RECT -2.500 -22.700 220.700 -21.300 ;
        RECT -3.500 -23.050 220.700 -22.700 ;
        RECT -3.500 -23.450 -2.900 -23.100 ;
        RECT -3.500 -24.300 -2.900 -24.050 ;
        RECT -2.500 -24.450 220.700 -23.050 ;
        RECT -3.500 -24.900 220.700 -24.450 ;
        RECT -3.500 -25.300 -2.900 -25.000 ;
        RECT -3.500 -26.200 -2.900 -25.900 ;
        RECT -2.500 -26.300 220.700 -24.900 ;
        RECT -3.500 -26.600 220.700 -26.300 ;
        RECT -3.500 -27.000 -2.900 -26.700 ;
        RECT -3.500 -27.900 -2.900 -27.600 ;
        RECT -2.500 -28.000 220.700 -26.600 ;
        RECT -3.500 -28.450 220.700 -28.000 ;
        RECT -3.500 -28.850 -2.900 -28.500 ;
        RECT -3.500 -29.700 -2.900 -29.450 ;
        RECT -2.500 -29.850 220.700 -28.450 ;
        RECT -3.500 -30.200 220.700 -29.850 ;
        RECT -3.500 -30.600 -2.900 -30.300 ;
        RECT -3.500 -31.500 -2.900 -31.200 ;
        RECT -2.500 -31.600 220.700 -30.200 ;
        RECT -3.500 -32.050 220.700 -31.600 ;
        RECT -3.500 -32.450 -2.900 -32.100 ;
        RECT -3.500 -33.300 -2.900 -33.050 ;
        RECT -2.500 -33.450 220.700 -32.050 ;
        RECT -3.500 -33.850 220.700 -33.450 ;
        RECT -3.500 -34.250 -2.900 -33.900 ;
        RECT -3.500 -35.100 -2.900 -34.850 ;
        RECT -2.500 -35.250 220.700 -33.850 ;
        RECT -3.500 -35.700 220.700 -35.250 ;
        RECT -3.500 -36.100 -2.900 -35.800 ;
        RECT -3.500 -37.000 -2.900 -36.700 ;
        RECT -2.500 -37.100 220.700 -35.700 ;
        RECT -3.500 -37.450 220.700 -37.100 ;
        RECT -3.500 -37.850 -2.900 -37.500 ;
        RECT -3.500 -38.700 -2.900 -38.450 ;
        RECT -2.500 -38.850 220.700 -37.450 ;
        RECT -3.500 -39.300 220.700 -38.850 ;
        RECT -3.500 -39.700 -2.900 -39.400 ;
        RECT -3.500 -40.600 -2.900 -40.300 ;
        RECT -2.500 -40.700 220.700 -39.300 ;
        RECT -3.500 -45.700 220.700 -40.700 ;
  END
END IMPACTSram
END LIBRARY

