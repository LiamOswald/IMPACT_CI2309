module BankWordDecoder(
input [9:0]sel,
output [1023:0]address,
);

assign address[0] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[1] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[2] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[3] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[4] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[5] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[6] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[7] = sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[8] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[9] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[10] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[11] = sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[12] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[13] = sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[14] = ~sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[15] = sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[16] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[17] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[18] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[19] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[20] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[21] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[22] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[23] = sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[24] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[25] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[26] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[27] = sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[28] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[29] = sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[30] = ~sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[31] = sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[32] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[33] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[34] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[35] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[36] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[37] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[38] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[39] = sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[40] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[41] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[42] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[43] = sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[44] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[45] = sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[46] = ~sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[47] = sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[48] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[49] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[50] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[51] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[52] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[53] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[54] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[55] = sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[56] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[57] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[58] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[59] = sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[60] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[61] = sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[62] = ~sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[63] = sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[64] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[65] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[66] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[67] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[68] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[69] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[70] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[71] = sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[72] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[73] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[74] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[75] = sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[76] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[77] = sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[78] = ~sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[79] = sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[80] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[81] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[82] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[83] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[84] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[85] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[86] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[87] = sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[88] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[89] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[90] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[91] = sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[92] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[93] = sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[94] = ~sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[95] = sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[96] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[97] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[98] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[99] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[100] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[101] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[102] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[103] = sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[104] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[105] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[106] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[107] = sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[108] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[109] = sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[110] = ~sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[111] = sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[112] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[113] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[114] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[115] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[116] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[117] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[118] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[119] = sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[120] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[121] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[122] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[123] = sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[124] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[125] = sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[126] = ~sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[127] = sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & ~sel[9];
assign address[128] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[129] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[130] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[131] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[132] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[133] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[134] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[135] = sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[136] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[137] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[138] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[139] = sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[140] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[141] = sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[142] = ~sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[143] = sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[144] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[145] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[146] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[147] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[148] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[149] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[150] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[151] = sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[152] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[153] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[154] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[155] = sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[156] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[157] = sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[158] = ~sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[159] = sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[160] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[161] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[162] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[163] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[164] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[165] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[166] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[167] = sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[168] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[169] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[170] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[171] = sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[172] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[173] = sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[174] = ~sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[175] = sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[176] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[177] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[178] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[179] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[180] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[181] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[182] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[183] = sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[184] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[185] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[186] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[187] = sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[188] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[189] = sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[190] = ~sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[191] = sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[192] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[193] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[194] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[195] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[196] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[197] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[198] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[199] = sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[200] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[201] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[202] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[203] = sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[204] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[205] = sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[206] = ~sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[207] = sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[208] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[209] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[210] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[211] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[212] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[213] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[214] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[215] = sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[216] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[217] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[218] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[219] = sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[220] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[221] = sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[222] = ~sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[223] = sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[224] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[225] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[226] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[227] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[228] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[229] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[230] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[231] = sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[232] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[233] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[234] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[235] = sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[236] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[237] = sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[238] = ~sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[239] = sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[240] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[241] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[242] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[243] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[244] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[245] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[246] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[247] = sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[248] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[249] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[250] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[251] = sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[252] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[253] = sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[254] = ~sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[255] = sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & ~sel[9];
assign address[256] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[257] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[258] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[259] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[260] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[261] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[262] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[263] = sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[264] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[265] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[266] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[267] = sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[268] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[269] = sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[270] = ~sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[271] = sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[272] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[273] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[274] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[275] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[276] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[277] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[278] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[279] = sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[280] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[281] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[282] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[283] = sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[284] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[285] = sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[286] = ~sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[287] = sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[288] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[289] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[290] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[291] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[292] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[293] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[294] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[295] = sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[296] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[297] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[298] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[299] = sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[300] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[301] = sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[302] = ~sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[303] = sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[304] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[305] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[306] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[307] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[308] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[309] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[310] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[311] = sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[312] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[313] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[314] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[315] = sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[316] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[317] = sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[318] = ~sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[319] = sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[320] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[321] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[322] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[323] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[324] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[325] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[326] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[327] = sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[328] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[329] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[330] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[331] = sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[332] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[333] = sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[334] = ~sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[335] = sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[336] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[337] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[338] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[339] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[340] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[341] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[342] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[343] = sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[344] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[345] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[346] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[347] = sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[348] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[349] = sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[350] = ~sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[351] = sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[352] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[353] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[354] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[355] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[356] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[357] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[358] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[359] = sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[360] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[361] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[362] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[363] = sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[364] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[365] = sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[366] = ~sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[367] = sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[368] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[369] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[370] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[371] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[372] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[373] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[374] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[375] = sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[376] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[377] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[378] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[379] = sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[380] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[381] = sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[382] = ~sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[383] = sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & ~sel[9];
assign address[384] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[385] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[386] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[387] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[388] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[389] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[390] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[391] = sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[392] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[393] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[394] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[395] = sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[396] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[397] = sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[398] = ~sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[399] = sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[400] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[401] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[402] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[403] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[404] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[405] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[406] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[407] = sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[408] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[409] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[410] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[411] = sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[412] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[413] = sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[414] = ~sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[415] = sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[416] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[417] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[418] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[419] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[420] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[421] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[422] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[423] = sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[424] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[425] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[426] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[427] = sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[428] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[429] = sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[430] = ~sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[431] = sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[432] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[433] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[434] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[435] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[436] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[437] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[438] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[439] = sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[440] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[441] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[442] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[443] = sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[444] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[445] = sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[446] = ~sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[447] = sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[448] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[449] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[450] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[451] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[452] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[453] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[454] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[455] = sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[456] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[457] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[458] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[459] = sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[460] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[461] = sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[462] = ~sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[463] = sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[464] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[465] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[466] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[467] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[468] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[469] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[470] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[471] = sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[472] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[473] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[474] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[475] = sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[476] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[477] = sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[478] = ~sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[479] = sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[480] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[481] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[482] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[483] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[484] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[485] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[486] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[487] = sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[488] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[489] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[490] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[491] = sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[492] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[493] = sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[494] = ~sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[495] = sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[496] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[497] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[498] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[499] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[500] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[501] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[502] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[503] = sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[504] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[505] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[506] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[507] = sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[508] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[509] = sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[510] = ~sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[511] = sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & ~sel[9];
assign address[512] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[513] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[514] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[515] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[516] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[517] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[518] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[519] = sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[520] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[521] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[522] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[523] = sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[524] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[525] = sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[526] = ~sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[527] = sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[528] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[529] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[530] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[531] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[532] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[533] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[534] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[535] = sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[536] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[537] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[538] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[539] = sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[540] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[541] = sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[542] = ~sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[543] = sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[544] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[545] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[546] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[547] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[548] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[549] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[550] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[551] = sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[552] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[553] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[554] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[555] = sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[556] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[557] = sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[558] = ~sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[559] = sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[560] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[561] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[562] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[563] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[564] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[565] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[566] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[567] = sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[568] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[569] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[570] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[571] = sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[572] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[573] = sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[574] = ~sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[575] = sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[576] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[577] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[578] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[579] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[580] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[581] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[582] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[583] = sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[584] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[585] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[586] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[587] = sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[588] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[589] = sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[590] = ~sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[591] = sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[592] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[593] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[594] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[595] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[596] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[597] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[598] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[599] = sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[600] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[601] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[602] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[603] = sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[604] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[605] = sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[606] = ~sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[607] = sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[608] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[609] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[610] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[611] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[612] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[613] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[614] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[615] = sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[616] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[617] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[618] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[619] = sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[620] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[621] = sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[622] = ~sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[623] = sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[624] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[625] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[626] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[627] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[628] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[629] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[630] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[631] = sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[632] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[633] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[634] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[635] = sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[636] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[637] = sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[638] = ~sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[639] = sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & ~sel[8] & sel[9];
assign address[640] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[641] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[642] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[643] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[644] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[645] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[646] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[647] = sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[648] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[649] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[650] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[651] = sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[652] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[653] = sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[654] = ~sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[655] = sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[656] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[657] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[658] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[659] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[660] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[661] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[662] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[663] = sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[664] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[665] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[666] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[667] = sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[668] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[669] = sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[670] = ~sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[671] = sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[672] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[673] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[674] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[675] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[676] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[677] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[678] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[679] = sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[680] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[681] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[682] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[683] = sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[684] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[685] = sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[686] = ~sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[687] = sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[688] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[689] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[690] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[691] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[692] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[693] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[694] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[695] = sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[696] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[697] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[698] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[699] = sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[700] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[701] = sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[702] = ~sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[703] = sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[704] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[705] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[706] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[707] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[708] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[709] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[710] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[711] = sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[712] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[713] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[714] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[715] = sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[716] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[717] = sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[718] = ~sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[719] = sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[720] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[721] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[722] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[723] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[724] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[725] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[726] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[727] = sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[728] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[729] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[730] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[731] = sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[732] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[733] = sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[734] = ~sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[735] = sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[736] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[737] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[738] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[739] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[740] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[741] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[742] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[743] = sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[744] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[745] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[746] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[747] = sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[748] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[749] = sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[750] = ~sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[751] = sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[752] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[753] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[754] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[755] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[756] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[757] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[758] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[759] = sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[760] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[761] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[762] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[763] = sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[764] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[765] = sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[766] = ~sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[767] = sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & ~sel[8] & sel[9];
assign address[768] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[769] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[770] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[771] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[772] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[773] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[774] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[775] = sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[776] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[777] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[778] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[779] = sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[780] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[781] = sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[782] = ~sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[783] = sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[784] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[785] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[786] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[787] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[788] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[789] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[790] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[791] = sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[792] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[793] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[794] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[795] = sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[796] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[797] = sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[798] = ~sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[799] = sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[800] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[801] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[802] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[803] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[804] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[805] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[806] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[807] = sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[808] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[809] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[810] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[811] = sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[812] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[813] = sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[814] = ~sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[815] = sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[816] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[817] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[818] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[819] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[820] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[821] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[822] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[823] = sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[824] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[825] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[826] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[827] = sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[828] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[829] = sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[830] = ~sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[831] = sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[832] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[833] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[834] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[835] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[836] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[837] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[838] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[839] = sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[840] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[841] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[842] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[843] = sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[844] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[845] = sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[846] = ~sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[847] = sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[848] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[849] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[850] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[851] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[852] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[853] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[854] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[855] = sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[856] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[857] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[858] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[859] = sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[860] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[861] = sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[862] = ~sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[863] = sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[864] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[865] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[866] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[867] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[868] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[869] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[870] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[871] = sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[872] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[873] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[874] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[875] = sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[876] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[877] = sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[878] = ~sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[879] = sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[880] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[881] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[882] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[883] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[884] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[885] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[886] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[887] = sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[888] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[889] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[890] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[891] = sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[892] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[893] = sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[894] = ~sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[895] = sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & ~sel[7] & sel[8] & sel[9];
assign address[896] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
assign address[897] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
assign address[898] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
assign address[899] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
assign address[900] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
assign address[901] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
assign address[902] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
assign address[903] = sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
assign address[904] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
assign address[905] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
assign address[906] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
assign address[907] = sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
assign address[908] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
assign address[909] = sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
assign address[910] = ~sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
assign address[911] = sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
assign address[912] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
assign address[913] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
assign address[914] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
assign address[915] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
assign address[916] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
assign address[917] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
assign address[918] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
assign address[919] = sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
assign address[920] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
assign address[921] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
assign address[922] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
assign address[923] = sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
assign address[924] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
assign address[925] = sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
assign address[926] = ~sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
assign address[927] = sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
assign address[928] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
assign address[929] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
assign address[930] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
assign address[931] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
assign address[932] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
assign address[933] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
assign address[934] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
assign address[935] = sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
assign address[936] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
assign address[937] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
assign address[938] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
assign address[939] = sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
assign address[940] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
assign address[941] = sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
assign address[942] = ~sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
assign address[943] = sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
assign address[944] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
assign address[945] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
assign address[946] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
assign address[947] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
assign address[948] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
assign address[949] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
assign address[950] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
assign address[951] = sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
assign address[952] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
assign address[953] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
assign address[954] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
assign address[955] = sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
assign address[956] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
assign address[957] = sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
assign address[958] = ~sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
assign address[959] = sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & ~sel[6] & sel[7] & sel[8] & sel[9];
assign address[960] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
assign address[961] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
assign address[962] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
assign address[963] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
assign address[964] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
assign address[965] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
assign address[966] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
assign address[967] = sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
assign address[968] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
assign address[969] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
assign address[970] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
assign address[971] = sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
assign address[972] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
assign address[973] = sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
assign address[974] = ~sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
assign address[975] = sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
assign address[976] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
assign address[977] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
assign address[978] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
assign address[979] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
assign address[980] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
assign address[981] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
assign address[982] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
assign address[983] = sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
assign address[984] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
assign address[985] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
assign address[986] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
assign address[987] = sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
assign address[988] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
assign address[989] = sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
assign address[990] = ~sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
assign address[991] = sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & ~sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
assign address[992] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
assign address[993] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
assign address[994] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
assign address[995] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
assign address[996] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
assign address[997] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
assign address[998] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
assign address[999] = sel[0] & sel[1] & sel[2] & ~sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
assign address[1000] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
assign address[1001] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
assign address[1002] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
assign address[1003] = sel[0] & sel[1] & ~sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
assign address[1004] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
assign address[1005] = sel[0] & ~sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
assign address[1006] = ~sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
assign address[1007] = sel[0] & sel[1] & sel[2] & sel[3] & ~sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
assign address[1008] = ~sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
assign address[1009] = sel[0] & ~sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
assign address[1010] = ~sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
assign address[1011] = sel[0] & sel[1] & ~sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
assign address[1012] = ~sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
assign address[1013] = sel[0] & ~sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
assign address[1014] = ~sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
assign address[1015] = sel[0] & sel[1] & sel[2] & ~sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
assign address[1016] = ~sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
assign address[1017] = sel[0] & ~sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
assign address[1018] = ~sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
assign address[1019] = sel[0] & sel[1] & ~sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
assign address[1020] = ~sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
assign address[1021] = sel[0] & ~sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
assign address[1022] = ~sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & sel[9];
assign address[1023] = sel[0] & sel[1] & sel[2] & sel[3] & sel[4] & sel[5] & sel[6] & sel[7] & sel[8] & sel[9];

endmodule
